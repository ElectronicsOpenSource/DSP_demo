XlxV65EB    85d2    18c0[�_`{�ѡ��8&��)��B6�`�����\�L��/�� h��KX�&���O���r�n�q?.<=�v�i�s�y���Ga��x��a�?�O"��\�O�4���kȑ����|>W��������	�F-z�U�K}�$I�+㘍��X=ߝ��Ĳ��O	Ă�?|�p[p_�����-�����|�CjvS�2qj��i��g��8/nC3S��L�P6.�|���Ѓ=�����,�큺����ż�2���6'r��O����0�HP.�m�aw��-eT�o^x���Ʊ���J<���lR��ۂ%Ò�j�ATG�����H�ȹ���c5M�?h!5�޵�?��.�G�1�%M�gK�;�W�
u�_��p��U���O\zB��>�PE�������XL;e9G�n�9칍�'�sĖ���vʹ�q����+Ee��a��Ҡ�X��4���؆H�r.����,��],�B��sQ�9{ybd�Þ���L�'~�1�a
�ZU�Ҍb*�
�h��O/�ָ)��o��4� �H�LfqCmVr�s\�%]q�c���Ш���ٶ�t��0"�%j��h�f�a�yw���C7�Mݤ�����2�r��~����@�!�`�p \X�>OoRM��c�n�C�~�idu�\� (�U�`�gڼ7btcwxΩE:X�ҶR�\�?{e��YO]��@�cL�q��">Ϭ�	��/�
���	Eq�}�9Pp���	T�~�>�U*�s�	��7+k��y8��ꮞ �m9���銖��[�W0�Ӝ;Vn7V.�nw7��m�h]O�wǵ������V��s���`]0���Ԇ1����j��Q�6�߈0��g)��w����8|2�D/�]X$WK]�o9�����ձ�z�6Aa��@1F��j$�9���j�϶\���=�n��L#�M�P�5B�z�QE���s������`a����(��o��������֮��U���<�!'�f6�0a�2���а�Qw�����T����S�d��C�ݿ��Q�@�u�)�LW�`{%8>� �����c���26 x2̜�K�ş�p����'�n��\��P��5�D4[9����@
=(=������j�Ź7��q}�v	l�x_�8OT�������13���{-Ol<f�̘����lMW^�~�ʷ�jy��5&G�Z+���-]�?y���whӌ3h-Uv���*~�c���DD_�Z��%���'[�FY�ݯ1 ԫ�����|�^�?/ϛ�('`�Lنy�y	���jN��H��W7�r��f��[U���Գ6�g�}n�7�� ;�* 0�6y�����^�@.�fIѸ�;�G[M��h7A�� c{�(�)9,~'��G2��6��k��ˢ"�{u��IT�1��'�՞��Z�Q7G�D��?����[v�������n�A)pgřl�B"��<��A'�0�;�"�]��u'��L��3q��s��Ny���a辀	9P�aq����N%�3~&&�@�S#ZWc��5Z���K�֌��)D|pgjI���m"D�;�UW�eѶj��Ud�-=fӪ���n��7�ܣU��j@�a䶀I��l��{T�f^�ƪ�}L��;��	�⍨q�=�uw�3;T�V��mU��nvF�75��^ϫ�a�k�;�/|A��[�����Eq㼔��%Zvp����矍~Ӿ4&踀�r=�L�`jQfA�z�Dչ�#"{���Ο�|���j%��dyeϴ׀��}�<*Kত'y1�oȃ.;s��Kmv�^_H~���x?�;��֓��4(`l']m#�����햘��޾i�UO�T�����Z�����6|��tc�C]p5�P���[is�n�`w�"��n�0��xj��U5PϦ�ݖ_+�h��b�(5�BYۼ_�:9n?����ln�(�>�!���F�j���B���kc���r�m�O�E|�t[�(Y�n�0LZIB�y%��x?��9ѤՏ�.؂�5 �;a��/�}Q�'T���3�e�B6�tel�T��!gm�)�	h����1���U�6��Ƥ��N�!'��cl�*�f�uE6@b�$w{�	@�{�Z�����ԅU߻�X���*\�1��˅G��]j��� _�4�>mj��8��X|_��e��`zUP��>���C_S2I\w�_3׼��6�t����^?�)7�6И.����3Um��4nB����C�4������@'�Vi�nc%[5O:��3%O��{�,X�8~���r�e�-�ѿ�R���md���,���#|�P�$���ƍV�CW)�x�,��L��?��ڥ����`.��ߔqE��G��gG}e�h+`�*п͆���7�����W�f,��ǟ
=��Yr��$%�(谖qX�ޙ�c�����S��ُ3 ���?��^4g�a��D��;�w22�g�%� R�\�A��r�
��g���Z�_Z�_Q��kB�X��a��=�!��.�>s	v�Q�<�g���;�^h��%�q�f������!���Yx�Y2��b6}��M-�dL�1s4� 3w���`�6�By�-׍��(B�rb�8E;�EC��|��l9�B&��E��P5��஛a�I�9܍hr-vJ˨�I���i�^�IӺh*<M���q�����6H�~�}N�H���4{{�A�q�Q ��褾��SY?>�!�v�WBF���^�E��n�Fp��*�~<R��$�	��s�l쏟h�"��U
��_u��^I�hٲ]�̽��X�=E��p�

�x���y��y�l�F@�r�*�3Ԫ��|;MQmԦ~�/�ˑ�֎.�Fa�;�.�o�S�.QG�[�WȲ�hc�j(���@�]MH�v���x�){� �{m��	yy��1��ك�'R7��.�+����c5�N��K�٧/��_q����7lT;}��5_-t�%*�G�Թ$8��k��9��Ӡ5�3��,�qj�w�k�V*�w��u��N|�Y�V��+��ouS�H����l��3�b��}k2�t4�s�6e��Jδo�7�Q��Өo5ˎ:�-� U!��D:N�ҥ>7*��>"ͪ�r���s<�Tv�ELmK�~3��zY�.6�h�!�[����Ǒ1�n�!�Y����r�[��6ы��<]�LJ�ɐ��F�=-Q��ʚp��)L�F�z#2��N8�M��n$�tK�eb]I�Cc�=7��V�	VxP����eiYb��߽O_�{te5�U���&�Ι`�#���
�3�LR��*�ސt	��s'K��U�,Wv}��tzZK.\�|�Cj\���vk��I�vƗ�Һ��/I9����e�_3{��=޳	'ܳ�j_�{���k�D�jo�\\�4	;�c8T���!������g���8���ɝ%�}\�E�+
��<>��㙚��;�Se]��)��-�}��������Èh�_,4�@�((�r�3`х�y��]�¬1P3���/��;P;*�Z��V�1�h�u����Yc$�O���O���b�D:����Ùr|�G����x���Zm��|��]����u�>l�i(�G�!�"�I��0}�E7��]���7���n.��\wȼ;{1V�&%�WSR^�Wq��^���8o�.��-��W����Ň4"���N���7$�� rا�17C���])�xI����J6(P9\�/S��1J�t�ji��N��	|�;�t޸2ޜ�"�U�oM%a�0�U'��a�+�)��g��u߫���ѿ�2���:�f��ѳ�2��� �<��|3Q~��p[tI�3�ê9v�b�s��Y�u#L�l;�vL�����_��M�J���F�#.��I�e.�_�ȵ0(�`�i7&a����or($ޮ8;���⋴si�ۗ��o��6�ݱDQC��hiwy��sAC��&>X��s��ƈ&Գ��pM�ɑ�����n��(�ߕ���O�p�-&���{ �)鵍d����%��RS⬴+�}+Y�v����0�3Cp�;=�Q�;�Ws0:%���F�J��ӴяaуY������W�+ɋu�����#�<Ύ%P&
�Ras�'��x����~���a�&z�_��q#�\�%�:r�H�^沌hOچ6�Y�S�_��Q6n���ٹ����W�IP���b]4޹�P�6���`ƚ����Vdku+�S�	��bn��� ��h���3�Y6kJ�Z��<���B��b) ׯP�lqϷ����&�P$q첪V�_���d���է.�OoŌ��ZLW��ۂ�XP�M"���\ޘR�f��-��g"�Ȁ�֯�����]�:9��eN�;�R��8�� ���P�b����ۡ�/�}[�����!=������_�r_���LO!ҍ}�T�%�J�}�-���+M��ڻ�0,3ͫ Y�=���ݥv�UoaTݠ�.��!��ݲ����a�I��I�\�6]�LJ�S�8�����ȩ$m�ߎV�OTM]�7`��O�����] j����h"*�
��G�s�8A����y����sp��;��P�8|_aC̺�0ذ� �!�Z�( #��/D���0oSy���c�����!P�t|��*�}�*9���3H�~V.�/7xOj67�o<��;�UȻ/k�Ȧ�祾~���-�sjE�Ņag,�M"���3SZ�q6:���*	T��S�r9K�Q>"��6���&�]����?"]U�/�c���Ib���,���/�$Č
io���q�2��VK'�����NqL�R����3'�6�(Y��aE6�*�M��SӾO�^���~�m����Ȫ.q;�/�u�@���fՌ
��.^�Y��(�w��tp�i�+Uy��Q�p���\�P�*@��k�ߚ:J��e�7�f��pQ�	�Y����x<É�|أC�ɜ�<T�;�p��!�_�(,���Jkb��P{�!�Po�DjA��h��ot1��k2j_�% %dv팃��RR�+��D��/0lz���\fP�����"�\��"���>%�;#��cȒ$Q/���<J�7��ocMw�0�з,��Y�k�g��O鐄v5.}�z�c���� /
>�9��>�u�^�߼֢☡�v�����5���d��"�I!~��m����u��F�����ް�N���,��J?�<rgݙ�ᾐpS�pvΩN߶L3Ժ�]רP�G�.�J� $	� �*�L�+�1=��<��)Mcgs\~Ϸ6z�M��W@��(�6��̫��Z�ހ`[d�LK��wb���!��}�$�<��\�P2�F岩{NXe@�J��d>��h-x�D�?h8֡�s�2����l?���Պ��L:uB:4PD�#�8�C���sS�먐�}64�-�����`��n1:Y{�n|s$e14�VE�K���t�`�1�n�nKl�ʽFt���ue�)�o�w���,z�� K���=�Tl���jf��\ ��$a3Z���z� ����?���Kaچ?�5�k��V�'�qQ�?�Aqz�	����ޭ�	o���3�×ReU`���8g#�PvV��
�~��Y�/Դυɝ�\���z���yh�x�V�g[�	O��x��ڳ�����(�8��{5�(�ǇN�7�����b��� �J��{�Zk풺�C��k�R�"�>5�ʿ����0�]�U��C���ڌ�w��C��z-�Ѹ����p]T�'83�%��L��x��g�Dn��8�8�j����3ƪ���^ܺ/�*�9rI<�"���J3��v�I(�i�~�� z-��G��Hod\?*d�����~�e9��T]�4��H{��2R��E���Oʟ3^)����+9�������S#do^��֥���l|]&��i���z�����&3�n0��"�}1aQŦ�P]��0W�m[�,b���
Ăx�5��EK��^��+��QwE׼��io�u|먚of��m�?t��ȸ�e]W����;�&u��{��NY��~�.7V�$��9e:٭i�7T䏔y�t��&3�E�S��{���̻���bw� �]$��(�w��/Cd�6�5b�}L�%�A+�4�ra��BŽK�*���Q��)���v�m��S�+	��ב|�f�V�s����)ⷼ6L5�n#��ɩ�f�@|vM���L���.�����f,<l��Rۼ��%�	.��ٴ�����UN���+cC�N	��{Ç;V�Z��F���Urƭ<7e9�@�����u�:�Ėf���p��?�8��K]�S��}��|�V&�
XlxV65EB    18d2     910�W_�O�hhh��J�#3��Y~����Y�+��h��^*^�uW���f�6���epL���@�
/��zIj�˵z�E89�
��%�i���W@;ows��&ysU�?�	ހ\d�.�xL6s\t�55 ����S}��������>�f�:����/�K�Z�V�*`�!z��]JT�
�A��)�R�HdN�ѣ���H�Ðfu�/����X�6S��.Er�JqS��nk�R>��Z<���A�$N��TL���ݳ�^�a\nܖ�nӪ[srW�n�ݤS��?�Пl�V�}��s}�3�7$��j~@�S����m'y�`1�� m���73�<��RR��@U�Tx����f2T�����%y�7 H�,��#��Ŧ�����慰C�}�Z2<G�1^fG�OJW5���=R� =��[����ɓŶ��]��J��J�_�bƭ�C�2?E����$��UZ2�?�%{qn8�+AO��]oM십T{Y�,��[C��\V�Vבb�h)���+#;��ꢷ��3�z�2�j�ƖJ;I�[s��������D��\v�Q����g��>��nI�G��g�N��SԄUu&GW�RR�s-Ӄ�R�۬n��X(pI�7��<"��u���:Z¼)�q��A��"�+�Y��Tm���N�3̞�^�9��[,t�t_㴘��:l
M�����)ŭ�� �{�V�v�/mL��+�����F�/}�NxF�>W�JU�bm��En#�m�8O�:�<x-�Y���?q�{��Qu`P���r��v�/΁��b|.�7_���}��f��{b�8A��h4�r�<�
g����c1!S�������J[h|S�>R\�y�NP�&�kV��-}z{����+z&
���F	���=�>�^0�֡�9�"]��8� ��Z݊��\�Rϑ��ziH~<	���xbL3-b�r�t9LE<ГI(�����4�� _B3����ո��ݏt��G��Ҵ��Jn�����������ٮ����A�*ȁ�Q?s��p��l�I?fbyG^����w�.��k_w�;<�v�C�]�����'�W/�=��C�9k�(�(�\'6����X��?�s_	G��'3H5ᖥ��Sj���`�i[X���,���|6G̖_�����k�}r�a^Qlt����`s���"i`���OV�/T�\�.��4�{�ٱ�ڂG��БG+�R̖Y�C���h|'���hڭ6o�U�=��jld NmB� �lzcG���Vʢ�(�nÁ~�^ ��u���qkjz�Q�fl���"����4��*d�u��sɻ���Y���l�;v><ӳ��@�nR��Pp�����ѕ���W&ȓ�# ]��]Կ�0)�<|�Q-����
UD+�)�|��3�B �FrvّlҰ�WыP`<��m�铍g��9�������|9T!��H�#\�����]���E���������]^@R3+���٣�=��qa�k��a�x�=|��f���@(@�oq��c��˲�;�=�K�Jk<��y�B�.��k�2�6]���@ڞ~������PٹT�����O|�q�.Vt��P���p����>���g���Mm%�SR6��f��H=�τ\��DD8�o#|�"�)���v�����*�ME'`�3�d�]��Ǫ��Ԛ����4m���x�g�a�7�j5���c����=w���Z��h/�&�3��	{>��1Hi=a���
�W����7�I �����֘�,D����*����4�JvT!-��.�D:h!8�e[Ď+7&�yfo�h�q	8�Xݵ�I&���,�üY�]�D��4G�@�IK�z���y�1ַ�D�Am.��ܰ��#�e����~t0n��_H��u$��"u�ɾ�6%���<�M��\��<��k���lX+�8���=�J���*�U:&�Or�1��O��II�� X��)v(B�}A�\:}ι��aU�TrJ@H����Dz4y��ܼq�]oJ$�c���f�y[���������/����/���ቇ_���Xx�ce��|���,A��)���yH��n�I������	� ����l�Ͽ�k��� ��i��EF��7���br�am���	yR���]�������E��U�����Ow���iJm{��f����Vy�Vrۚ��H܊�AN^ku��`��ڞ�9g�	���������v93��|��,��dF���Iޖ�/1�9�Vg
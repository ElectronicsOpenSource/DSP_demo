XlxV65EB    40fe     ed0��b�VI}�8�
-"�٢|*y�v8�<�m�a�I�˕��Ybm� �#�%��BHT�Ǌ����W-���~��VUn�̿��!�6]���Ef`.���Ј���H�^���W�G�K{���2�*�R�6�A�v��:�WhCZ7��J��B+,�����Q��H���!;��]����.2g�Ax���A�"�1C!�}"�tF��.���{��"A'x�R6hI���.�#�b2�0q �;,JkR��KChe����7N��
7(d��t[�P #uN���e��������,���M��&p[g��;0xu�ԕ��g��v�cM��i�l< �d�,'O�#�Q�HM���%m+t�����|�kR�Oc?bEs��E"��O�1�ۦ��ӕb)�j�vT��, � �z��uU��-�y��Ma���
p³�� ��pB�Q�gv�_q:+����Đ/+�&��i�Y��ݡ��\�VԴ�P����뀱�3��Q_�~񢱲��1+-!���|���X�E3�cb%�E�4���6�<۽��rh#��v)��eK�}�$}�+���Ќ���K{>��w�z�U�q�;'R:s���z��� <}:��/,*Ә�?��<q�L�� �0Gv:驳�3JC��BY���U쬰�c�^A�dI}�'�b���;��i��]�p�Ĉ=Ɉ1���m
@��1sN�s��ت�@f�x=�޳���+wXh���ȸ̧_7�
.�������?�+�Й
�.y=T*&ߓV�4k�,���&<�7�`�y>_�K=����;�ϐ��**���r���T���N��w0����;B�l�+��A�f�A[fl$V.?>��_���T!Pl�қةh������eL�5+�[���(�ؖ���8��0`�}$��j�=*|���Ă�<_(�,b�k�+#���{���o��Z>�M�m�oY��}��h�!��J�9��X�}��= �J�H�k�H���D�\/�/�D�x@bp��]���vM��n���;R����-��� ���Q���j�Qϻ����0S��)(�5�*9zd��A]�8�N�����$�y�)o!;�7ÉF�����/8��;��#�8��I5�3��m�NuY
���&�$lZE��$
�ƿ?=�~/�� ��7�)a���8��:yC+�땙�0g�9+%Ah�hő����̱��ws��Ć�8�"�kA�/��zf����}[���(D=���E�.�
�
�lH؋��t�ӝ���d�>f�_(uV����>�f�@��<�fbO�/{1[�����;����AK0�%_X��Y���Q�vDѶ�� &?���^� '`�5�W�J�Gw�3��	9�&Gi��3�\'Փ<���V��<5/o!Į�_U�GH��E5C��Bx�џ9��	�s~�<
�Jٍ�|5�xC�x�<C��~���Y�iǔ寯c�حT7�|���;}7��7F;�/����I��q���JB�4�N[9��"Ԣ_!�����|�#�CE�1z1?Z�x��o�gӉq�j(C��e��9�B�"�z<�Ȧ쨊H��T���X��M*V��)���ic��|}��!��0JTGW��s�8�`��'k�ͣ̉Fg�^j1R֐T�Z��wi��Vy����`kZ^aB����bϹ��ҝu{
1�͘����:x�&u.�݈���Ғk�m���ղ��Z�8]�������7����ˁ*o�,��Kn�������Ӕ�VC�^r�s}�Y�}�C���=�6S�N`{9�e�C��9�a�� MZǕfޫ+;�]��̊ ���u6�D��6��0�b��Y�`�0	��L�햒�\�f��v�_�6p�Tc��k���9�-�D_90�]�3Ii��we���+pd���w/��F���^-5������C�x�4�9�Ђ�m�өP�wz�nlY�N‏�����P:>�(-��$W���=��AڠAJ�"�ң��м�q��T���!�]8��2[�7����NU\����}���ʧG�WO�k�QT��k~ie^�q����c��'f�6_�InR�:�!���d6L8��h-ӊ@z���nf*�ͳ��e�����c�_�����,���c�h�:j�䓟Y��t̐"�?/��!?��(9>T�1��s�A��)?���n
hT*���3Z�A�2�ah�	p�&��/�'y}g���7�� ��Kr��ݭ ��}L{�k]���(H�p\��C�@ڍAE�q���V);�gݶQ��E�)g��2+�B�9�0f�?��BWz�~��C&�"@�ιWۅ�RZO��s��)4��b%$��V5�\ת\���`z!���S�\��|oP�mxO]�
�e�C��2�]m��x+�f0oK�y�4��W�Di\��=�~�� �ӿ����S�W�~$q��h��]�!����j����Z�2F�Q�	d7��.gި�a+$�B��&��L#ﺐקv��ر���ͱ(��f9�J>��|u�Gx�	۶�8�E>�������|$\�M	&�z���G���R��
q�|OI�� V�<���8�M�\�q4�6	���3N�ed�^b �G�&=G�Q&G��^��^U�i�|%K&h�\c4L~�7Q|����,z��3LU@��6*O��v���mgd���&ǂ��ݤq��a��|����/_X_���u�x��!��E����F)#��u\j��<J��:s��nE�
���j�k���ey[/��t���yD�����]c�o,��U��'UQ�rQj�A՗�����R���4T�^��"l1��N46��G��ɬa����i|d7���e,�C����ѫM�Pqܖ�5����,'�d��u^�s���;B.6���W���"��w��!����"su��[j���b���e�ɗ��Ʀ���v/�<ء�
[�Wg�!�~K�&�?�4�e���(`c���m=����mF�)*�=�����0[l8S���ܙ�-���W4]�ы�{���TׅH��QA'Mu�S9N0S�E�P���][Gbq �h�=�ތ�|�@�l��G���܃��0��8�����e*b���  �o������ނzܢ����9�31}�`��P^�q*7���5#��Y��+�wY�j��`����P��sm6Q�kLfn��H��w�U�N!��S�l�%���H#�h����-[(�괧�1��tv�I|��҅�PT��}=�Ɲ9��§�˽�Ji�~�/��!�X�-i��r�ϔ�6Қ��VF� �����c`$ݹWZ��Ѵ�IY�HXk���ўd<��lM_TPl=�d�ق�
�@k��4�+�l�F��ݩo�����KS��
#3^��Ԋ��@O�hzI8��P�g��z�+׶&/��4:D�e��df��-'�N�XeTh�����
����֚�:E`�$2?+�`^��*g�n�C7�->;g�~">�Ѭ���'G)��lpb�6U�Qu�R�	z�)�l��NL�m��D�1�2�q7�����D��?�Z[X�tYKP�q�7���mCB�U�~���=|^c��ߊ�P�Dy[�{�"�H�N�^��B�w�W`nSטl�����޴����CF�z3]0�ۯ�/�\`<�^�]�d����@�g�:���i G�Ak.�`��: �O���D��JcX.��o�ݳ�:�� �D
XlxV65EB    1f58     ae0�Ql��A�=��_b=��������c����(ў��q�(�ka�G����F��-}�df�_O��լ��Ke�&�[/c�JJسw���uN~`n�
��izu&�Na^�h�Ra��p@�;M��[��E�?fG�� $�8�z���1���(\q�:��%�����c~<c� H����J4�5�--E�Gz��p4��_(������ACk��ӪH�7�ףq�~j1�������Bq�U7B�u@UJz����`ǂ�0ϧ��רI��~�oI]p���M�'B��ro�����a醬	�����D���{�[;-���@/z�j|�w�@y�pg���NT�vG� �YjJY�7$8�s	H1�!�����d��=��d'Rd�S�n���\Z	[��7T#��c�V�f�3��ֹ�^��%Z(�� ��Ÿ��c��9�C�l��(F����6��j��	����wB�.���wZ�����#�D<�~��.o�_]v����@�IW�z@T�(z�_k,"1�:;��/[��`�߰d���2�*M�9W�σ�Hi$�[����L/>q��-�H����(Y����S˾�k�.�]O8�Zc�Ez���Ƈ�=�Du��}�	��?b��k�R�JQy§�@��_:�we����ʳZ�k^�/�_�S�0[x���U�&^	�r�L�˞g|'�I8fU:�� �i�����cCT�o���M �h�PQ�d��Pr��b�e�����
��� ��z�n��7�%CY�^��#n�$�(��h�
��F� ��R}�g�cxd>f���q�:%G'��*��s8)�~�0GoS��5P���;?&��6ϐ^I��\��f+�����Va�|n��vch���)��1�%8��{Bj�C���EB~����v3J�#{�'-��1�TY7����V�m���p�w��?n;M{�¹�$5�T�"0�HN!�
��D���>dq)�X�}��'M#r��Е����_9�䈇��\���G�s��3P�p����T�D���us�Hfc3>�o7M�m�>�]B'%����{h��A3��cZ���8͏г��;���'��KmPN�h�G��m��|�'�S��]�6iΞZ?p%ET��;�O0�u�K��;*��s��¿�Ε1�Oy���B��v�/�N(������r#1��bc�(��[ϥh������4��?��F��RB��	��;U@�\��S��7O���KB��I8"Fo�� ���d��I��;HbxbL��S��W�#ў:!�v�:2������}��K�=�-�Jj��-S��E����ʻ�K/V�f���ۋ4&˟c� {yvY�W�s�DBoƭ��'Xb�Jh��U�N/;�r��f��Z.���^��>�����l��ג=�4�8Zf���m�n�O�(p�}[��W�]��Ԃ���:=0jp����G�1 1�i�S���o�y�7/������gp����pxn������[?����|��W��U��W�*�����~�,�a�zi0��ߩfU���J�:��:Ui{��D��G?�l�����f��kr�o:�;r����@\���o����o���"x��EL�)+j[Q�7G7���b�%�y�����aG�$$��)��R]IM9����i9ԫIa������Y�M�S�9�ۆ�T�9��y�*4�8�B���Ô���&(�7jS�:��̽O3��F�c�	���>ek q2��Bы��'�`�Cdq�h�V�.f�a�'�!���qp[���p���c�w)Zw�#ʓ:�i�e�&�^��&7�� �1�E���\�LH��Av�D�f�đ��y8&�&�j��Gmd��Q[.f�`mm.����wM8s���M�B&���&X�����Q�F>�+٢����rC�U0��C�2�� ��$���������3�<psr6,u?���h������X�g����ERFF�	���kL!p����^���>sG�k��k6�Uq�Ev�>��1'�X����L�W�F��u��<����QO{�{
���BDf�5��-	��ʋ�v"� �8N �H`t�V�]m�'=��G%�Ѝ�T|?�����6E0�d|6i����Ȝ����d�a���M��� �Q\�����<������҃H�=����v�-��]�R�P2�!`�?8t;��R_��U���&>8���F�-�!C5����!KQ�V�ھ�x��X���zNڇ��yrU�y�3�4��1[�턾k��J�g��w"��}ػ�t��S�9���W:��(. ��
�������p��p{�;#�E)�zQ�j�_8��"5�("`����l1�����Rv[XƆ�~)�_�=���]���>dD�7� ��~������#�C��E��	;���k�uvZ��
lĹ�t�50�zt8fW��Hƕ�������K���|L��z�v����9�-�	���Z;�8o�J8]m�~�u��ϙ
v,"8I�W]�����A�Ds���x	#QL�l�DW rUo�(�t���XdU�8h������ wjۉ��P��*W��|%���L������Hd|cqG�3�%�]�ȯ՘��B���>��'go��/m��T�*l�Dz^��*Q��{�u8���C�����q�����{N.�\�:�q�/��޼T`���c�а�}��Ԋ�L�����/zX��>����ͦ���:�{�� 4��R7=��
XlxV65EB    185c     8f0��;��f_j:V��)=q �/�9���M]Rт���d�AM==���Z"j�мA>���~u-��!GI7�����s]���/\,p�w�j�3%A��Ӣ����R
�&����Ҳ!.�E��m�� ��/�a�5	]%1��A���v�V9�@ʊӺ�]LFn#����L��!�ܷAĲ
�U�ȳ����Du�)�͛׎.dF�V�K�?��P�˅��E�5}�}��=�
p�4�e;�.؟��������m�˂|'x�/����R�T��K+*>����lj?���wJjh�֔^�O��d�/B�a�`k+M�E�v��_LЁ��IݗT�R☈%�mW`
�����Z�,|uO����M��l��d��m����qR3գ�]v�CHo;I1������/�ꞙ�#�BU�S�#/�i���;<���)�W�����.���D������S�)[�ԝ�`���� آ�q�AK�7b�׷D!Gu�ˎF̴��)�9����g^>F1eZ��!�K�b߷`�21���;kYܓ�rF좔P)|)�=��3�I���/�Qo/5|v��_D��O�3�[�9���7ו�H��J�f��[�ѻiH-��wI������>�L^�b�u�"��ӧ���{��Ў3���p�����X/)%M�1��v�@d��%H��.;}TB��|��``$$�F�4K�@S�W�F��Z�����U�����x��o^�:��$4�Juu�mu�ܝ�Q1Ĝ��*b�Gۿ��_u�C]C�yZf�y�P�!��<�#����˳�0��9T1�ޛcc��f���E��������e��m���]�3�	f�^w���Є7�ScȋU{���]���Z�NNM����7d���ojp34!7�k������3��2�L7���"���8�$Ei:Pe3N�g-{b�z[<z�aqG}��?r��;���/D�r�ߓ����5jxEu��)�L��ٮi�*q��O�g���8sMu�cF�B�z����KĴ��v���à،wu;XFӲ
[�����[qz��%1�e�ts&o�Eo����5
�Y�A� ��F���C�z}��������m�u��p��Y*��J_5�ɳ<	��qmu��8o�)%����c�	�\	�<!
p�d�'F�
H���	u�;�}K)+�.%S�A�7I<%��i�ٷ�4�*@��a�q��(��qgܽzެ{� �T� ���^�s�-�3-���E�X�lf��X6�8���bL��zc哭�����h��h����|gx�L��_������������c���ȅ���)�4򬆩��v�X�Z+CjP;g�C�l�	�FL�g�Ƿ���#T,��&��`s�$��`�c�0]ux-��4�Y�&5��Y� \��n(�`8�bNu��S4�����d�(����GUm��Zq�Y�B)���"!CG�=�a�#�u}��i$q��N�h�E��T|�|�1rB��7�@'~a������₋s��1�\���P�P��X1i��
�q�w��n�e���}rvŗoJ�#9..$0P��K�J��x�#�yi�fsPЦ������)�T����dCMW�3�M�Áբ^e�sW{gȒ��~��'�������C�@�Z!M݂?��y���"�F�Q�[2�#Tj�w��:%~00p�c�9y��+�U�9g��$� Z��{[	����Q��,�S�T�J�Rd;�"h�_���E�����5M�PXs�qג�~�ٹD|{KS�im�!3p���ly���Rm�f����FS��4З���v��۞�Ms�FI�ü�2;��0���k��I��J �!�\C^�#��,P�E͙o��!_3u��a�gv�zmlW����+�sG{��P�Ⱦ���=�3�!'�����o�?/F9҉}1��e���e$h�a�K������WkHGW��Rq��4���n���֬���AA�S�k�nș0Ɛe�9�	�AR����\/��u��O��֔R
{��4�i	56���9NP�lX���Z����*�h�iaZ��H�η������7ND�}y#�\]�:�H���Gh���������0n�ل�j�
��t�Q,ާ���g7N��2V� �
zxSج��N�R��e ;��v1 ��BW���R?���ו��y�g/.i4�^���Ζ��ޡ���ѻ�Y��a�(#�,��3bm�C+G`r��!d�'��?��.�N�-���eb
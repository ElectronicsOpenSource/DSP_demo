XlxV65EB    fa00    2ef0=�,�g�f�B���Ga$w�L���o���]S��[��eS�+�~��a.Ή6���tqI{�VCV`��'���C�I�.�a��B�[W���W��,!rg�=S~en�����$|m�j٣\�e �ʣ.y�8�ih�S����Cۭ��9���Oh�6닝شF�	c:�?Q�
8�t(:B?���Yib���A�EN���tZp78�B!M$����cG�#��	��i�*XB7���Ӵ�a� ���|/h����q.�[���]������@��3�K�^�K�����p�P�ã��Qf�Ғ��ː,MwYlM��,v�^�~Td��wHp�a�v~P����c���1� ���}a��Z�E�#Fެ�ah��0^9���?SU�"�+���'i�|I�<��N��rl[wx��ttt�h�󳜈���O?Ô���ཝ��Љ�#j&A��1��(Rf�&��*,�F6�f�k��P�Y���);ïb��L�C��
[��ܣX(��iw�dV�κ�xB�F�5�J�j���ܸ�oЩ�����+w�Jc���ySisj9�~���7��Oy^�^�QQ0� _w\l*�Y*?��y�wv��5������"Gm`Ǣ�7Fm���B��#�Ԝ`�2C\��Q�c�	S��c�	����}5.!�t�59��^\R�p�%���zosrgڂ<@^�ӏI ��]�<���<�����`�"(Z5�<�!��!Ò���{µX4�EfȆ����H�� �vs��_F!��pڛ�~��A�P�X��_����f/�w4˭b��0��)��c�)��I�Q�Ĵ�T��32��Q ��l!\H�01�w4޼N �>�o��ʢ�dM C6��Y9�
��^�'冀��w!�a9в��u���F`�� �o���M(�0ڥT��'�wPo�t�n�`ѩ!�v���������bՁ�޵��(�|q9���	ya7�����#�?��o�ߋ���1���a�8���p�?���r�����(R/!�����^��8�w�q�Z�"l�l�ǲ��m�?���e�(��^��ށO#�!��go�	�K��w�}�|��]k3������ �8��=�U�b����#}�1nb�8)�����s�V��b�-Xee#��I{��<�1ߺTc$���l�wC����D_~��d�z���r��b9f�5�g8؛l�Mz-E}���a�YaQ����bG^�}��]����8[J�.���j�ȯ�y���n�8��s��?��gˍWS�E��l���V���cM�BPH˗Yq��XV8Ԇ~'�n��@��m����ݒjA�_]��A3 �K�K��fJѠ ���-.U��u�<7o�:���4KvV�P#��9�#��R��&l�<5Z)Y���7��8��i7�$���6x������Q�8�q�n���~���ཙ�$y{�JE��Lt �꨹`���Ğ� =6�;X"�� B��Q�F����62�͗�H�:i�|ϸ����ӝ��KRF��ӗ7��d����V�����i-_�@飛��)�hYa$R�o����0�: �9�e�=�xg�{�tN��(R���tcq��e�Y}����k��.����Π�����T����faD�`Yu3&֤=��e`�%8��|c�GLX,�F�%�g�Oމ_���p��vf�K�zyM
%~����)����]'<j�2��ׁ.�L;iY�Rc�Ǝ�F1���������SF+)�zW <I��1z�5Ӵ���6*�<�k�u�B�5)V❉�]�>c�wM�z)�� �(
� E,�M]|GO��  n�T���L.}@�	s�����cM��eM0s�M�����f�1�r��InTB����eh	έ�ѕ��ċ5���N�z�]��Nln�34�$b��l�@p���u��w}�[%f�V�������D.1o��^P���ea�]t
�쇭1x����_aQ��g��Ԛ���s�`��@�a��q5�Zo�~����@gĠ0j��oL�����w�����<*��R�+�ƴ��*�� �R�\՝�������5��,��;�D�q�z"�Z��F,�CqP��n ^V@K� ��Äa�˰Z7z6�4�Vh�hBy�1�LE?k�&�m���볞f~��P>�k����u�2�+l��b�:����O%����8N���(�T�0�A��׿�5W'\�{�j%u]@�㥌�����Yn[oU���Su��������4<^�Eh�2��Ҳ�f	&/s�CMƞQ9;n��(��;�l��|'�����U�Щ,c�t7'ׯ�^$�Ƈ�J��3|�	���P�b��ǠKZ����]�՗��n�:V� ��1{lOݹT{�"F�l�]�h�%�YP�����Or̺�iC�4��hN�<Wrʵ{��@^�])��p�<0Y�T�D�-�9�j��})�e�V�t��7��FY�\�V%��h�߇��0lAI��Gb�.�\�� �����YIpJ!�<��s���2>$|.{�{��(�1��(���uL�!���yBv�l�@
W;�8l�˖}QWl��:ϚWh�ֽ~ǅ	�Dy��<�!(�B�m3Ċ��W-)w�ʊ2Q�ޕ����cm}�58��;*&�RS�*H����i��<��[���v`�7��-���>�G�Ѭ�^16�^%O��?|�"�Ɍ:h*J]�z��N,����H":��/"�~�@*c�ث�p��ʤ��ZE7��Й^��n�����R�UhE�m��rr�4��/J�."�����RM��Ws��x̙|˅�����ϔ:K���;Q�.�~�m�f�[�s䬒� t�{m��gE�:k+�ȑ��g/�<_S���6Y�R�F+����@z�����^��$M�'"@g�nI�r#��,��M��R)bb���fw����f��=.�g��(�k8Q�7�~�/Ҽr����)�(�>~�G�*������P�UӬf\���E�ց�@�<Y\X��т��:�A(ޱ�Aڧ�u������y,���&yJ,��5n�R)�r,YW������{ژX����)"XK`�9Wʷ݄����]lg6)	y6Lf.�j$��r8f׏��1�u�M Ѱ�ɫ��q��|�����K�*�x${��$�b�F��8^t��̿J���/��k�N!����,<7�t$kZ�MɁ�=�6����4L�PDH���v^QI�6���F�ϕ	���^r�7f]ָUV��O�~��QɈ�f�Y�L�ZV	�߷�1����sS�c�8��'no�D�m���J�
Ɩ@��uG�EA��.��
{��}N2�<���d4�e:k�P�!Y@K��Ts>�� r�v��i*٧x$��95 a�ق|�y/��������z�@e���m��N��2�&�7)3�4�ւ8ˎ�U����8j
V�k��齝-Vz${�̚�2�B�/�\�#T@��죲e]w��0���/u��е�猞�`<���6�:�f�a�`��*�z<��"���ߎ�.{UGy�?�WGO����$yc��l��`R5���:�I��G�km���v���ۗƜ��a��o���D�ri�f�r�f���K �䞤�=(J9��8��5T_���S�v��āM+���!V=団6��2�� b��;hE��x:�Tuը�A���on{Y=��GSg����*�E�$�C��'��{����g��qW+�f�Q&�>��K����'�S�,�-*&v!�&��i�7&^[ns(T���	�$�0�G���Y�Z'V£K5\b���25b�?9�Ȟ��q��c�Й�Hr��I�j�s�v^[��q�4�ۀI\��c�lӊ��}��4l��`X<ޒ�;9�>������]���*ك�e�dF�=���cZ�ڛ�V$�?�~9f�!D�+��Mb��8��!���T=��Z���e�<�&-�ak2"�X�q�6���S�"2��FX���ot�l�ɼ��(�BR���횈�!�>�!����"���֯$�"�[��t���n�'��r�-���/�(<�bb_��q�By�SK��'`	~��.qp�U����E�'Q�N�����[G~�xQC����.]He
l��\��{����1Gq:����=�uUWXڄHi$(ʪ����1Xs���ti~Z!�DF��H�z5Fv�M⪸�/��
�n��B�iD�})��A�e�meS���5��&?��F�
1�=��e �H��r��*dıJ��<Ԕ7�dь���#�/���!��U8�!�Yx�쿐q̀���������	��!�ЩD��/����KI��'B���s����Mt�g,�V#�>
���(�PU�VJ Jhp�2�g���h���r|�>N�኉�㑡�k@T����� ���<M ��b��k�r(u'�� ���eD��*��x�hW�ټ�%n�M�= 
��@W��upq��׊N8�f0���^2�nl��z�B&�,�]u2ا�3P�Dm�X�����ǽ���5R�v'��t�i������1-@���G��U���5z���P'�R�����'� ѕ?��漓h@2<Cr�BG؃���{�����D�hH*x��xh_H5���@�e\��.��5�p���� �Z6�XR)>���<��E�x�:�w'$�ގ*�w�h�|�Y�U���͖d�Q����u�� �� �Ǣ�t1�_,�Ka��{)�e���
�_W�m�H�C�~*(���M�/ F�;[���צjC}Ɏ�����D	YҮ�/�@r:<��P��̃N���xC8X�s6Y��}D���08A�y��#;i C��iF�CHp<=����]��4��7��N"�H÷�fr��l6�:�~<��3t����X�HOp:�RQ8��^����Q�d`S�.t)��,2b�����ӌyum3R�o);˂ 3̶M��m���d*�,^|�zX�ϰ�S�Gs�z0�6���ԧB��^�p>H5��[���N!O��kj�X[+�̶���v��eU)sǸ�<��ϯe�J ?;��|��IC^TX��x�,MFr}p�ކ�y�!,U$�V���~����K�^��?8Ca�X�fk�E�hs��;~L�rޟZ���ٙz����O*��JZ|L0l�;����cݰPƄ�����x�	q�I��M?�9���s�E�~&�> �KL}P��'�֮�QH�*?���Vp����O�&�)�3��j�˪�6�N�!�0�U�A��<8�;Z"{�֏��D�w�ⶲ�Z�uK^>Tg�J�߽�O���{M0
�o�9�܅��]���� 5E�
��;EUwDI�$�w�Q��Ҍ����Ud���[�\��c��
�䎖8�kt<P ���&J�����5��x�q�+��2��i�8'�PT�^+s5 b�F�
��N�vӷ
o,��R��h����:sCf󋎅a����^ ��ԯ��Q]�-����˰�/ݹ<�c[���ǆ���_@��Қ>q,?�#�׮@�	$R�=T�\rM��=�]��i�g&� D�4� �*�lTˍ�F�s>a���6E�.�Ҳ�e���?�'�(1ShYdM9;�1i�l�!�O	�y����t��hh�c��쎸��m����;���F�]��C�K�%\� �%��=��H�p��g�Q_4����A�x�O��P\SK9�������Q70�f�������Ar�:�*����w�h���Si�P	W�q3h�|���
�Y5���M�H��F�U��E���)�ޒ��e�=���v䊊�V��"cL3Ѵ�.��V{�n^n��G�G]77��<$��<Bo��9m[�5N{3��4��,���t9������5;]���˧Č45���,��I��'K^֌�(���8���m���+c�L*�SK�5c�)	_��|��o�ߙJ�ˈs��?&y?�:�0q�3l���1,���vՐ�b�5�2�O<����g�[Eg�6�$��9�d��`o��Zq�_9,�YnʱK��hN�Vq�ϝ����Ns-�_^���pK��٤�2P�D�o�$�T=@!{#�ȃ�Z�ga%Vď�
0!ե݉��jLf�d������3S��?��"�N�<?�����x�ԞUH�^�	É����e�0kq��� �������n\���2;��Ƈ�0�3(i�PG Ʌ�/@�D�!��z�ྭ�[�4��k�ڳ��K��w��,Bco���?��wP&�)����u~t�#�p
��)�;�0.W�9��y�G����(�1�ŧIzO�d�9-	|b�hc����>+˳�.�CվJ��Q���F�7��t�̕�w�7����Q�E�0��HՁN��9�6�\ RV��᱐t� ԕ]�Db�\��8��=�Q>߷?+�?#��3���䬮��_�.���-��R�;3�8HW�z!�@u{g؎���3�h��,z��|_���),}�mD�u��7����ʎ���̆��;_�/�9J�����t�;3���}j,HoWf�!��q�?���bl���*��@�JɿM�R6��K:数��(�I:�x�a�%%�2�%�Eͽ��o�����{V /�H��Fu�k:߈�#k��M�[	8J(�3����y��2v돢��/�W#����9�ꟸ��c�-�&a>��č��?�4N�7z�|���Z6��֠]�;��W����"au���j�Ŋ9�O�U�ZO��]�&_q�V���f-T'����'��xU���ф[;�C��P��@�Lgȇ͚�i��B���Z���P� ߀x�vB\���K1���oXoâ�6�P2�1䮽��Wt�STQ؃NY42]$��J��ĔWPqo=!$L���?y�v��~T�9��[�	��>�fo�^�R"�*�mB�}v���%,Y:R��6�QYJ��Ӑ����u�?�5��o:�5Un�2�K�&��	b:9�!Ȟ�]��������y�!_��L�>�z��r��6��AF��W����(��s ��y�D��@���Ea?���TRq*�({d �8��秞(���W3e�GS�.\QJ��S�pCLw��{�w�I�S=���ך)���\#�j52?=UVI��lق:�ЍݳMt�g�Ѷ��	u�'t��)���1Ϋ*_�-���u�>�~�RH�����X����d���+_Vx�@[D�i�[7F�*u��u�ˮ�t`�<�y@����t!���Y����#ǳ�����vTǓJ���E%?����Q����N����D ���c�0����8k}����K�GD[",	���3�D�M8�����9�jS��R��ػ���������Ij�M Ҧ�f�!V���ѳ8p)��J �"��st�O>��)ȫ�mgӌm*L�XQ�S�Cl]@�r�,�q����[\�G�d��r�~�	�Y�!*< ���mw��
h����ah4�+�%�,�*a��h!%5F����i�U��;�|�s'�������#:%�j{n���2z�.�i�i����9��Z�D��ư:��1�,s@y�2d�H�o5��]���8:꺨 �~MC%����?h�i��',,��,�z����.!Iޞ_�g7p�!Ͼ�Bg�����i��I�Y�Tk`��	m�[�m|�i��*o��r�-p�bp��P������3�l��l �~�<v�}lf��/�bѤ�I�$���9^�V��FC7~3���]�~��77@�ީG��UI�p^͸�~��
�~��+w~�4�|}���q�����9�:�ߎI�zlC��Ha*uoҁŮԿ��#���hvg۴�����Y4�q�!��7N;�/�Z��~zŪG)j �ڡ;�W#ʈ?-�^�LL��L�T⟆��{����c-���;�, �E!+�^�K
&���,K��k�mJ|�R��ze���P��7�����)�N����<g��Q�����|��l��L����|����+���Q%췷���]}.��h��'��c~���~_�����p�9X=�}-�_�HX��R�W.f
b~L�������fQ�w,�2�H5� >�#C9�^SO�x�)yd�Vf#�G�}k 
C#q嫿��p���Z7�������'q��QN(���<��*Sю	JCR�}LGK1��d�S�����F1f���쯋ֲp�GXJ'��&�\�T�Itm���޷Ҥ�|����*��T~��m�8L�WC��8F����`�cR��b.��W�Jx����d�$�JMKVن�Xe#�v��k����#��v��у���M�)"���R�á�l��_�)$�ֵ]���p����X�b*�u�B�dBc_� �ɦ0�OC;+��b�%��� �.B��D>H!�R�.B2s}{����	0��9C�������-H�9J��0�X!�K�@�p�GUC.Yo�%���V�]�j���H���x7�ɲ�˽؅X4�O�J,��y�ޓ�'�l�/!�����~Ds�VZ��%��W���.e�l�0�7ǭ'�U�mJH�b��0qB�u�?�5��P���2۳km��a:?���,����SW)��ԏR�=�}D~C@?�|KW�v4r-NY��WR�j�2wZl("P��@��(��[��\ڪ ���T_a|%��*9��"�J:fh�-��la�~�HV:�r����o3t&К0��
j:�;��,��ĜI� ]M�3��!3�'GS(�W�I�fʖ+ʯ����O��Ӧ�s,7C��A�6�خŞm�8��+1�ʆ������5�2*&���&?p�Y:=[^>pR¤�ϖ̗c���#��w3w�juA��.����*���|��i�G/◥�9����l�Ԃi o��Hy�IU!�&��d7�N&���"�,�P���Dj���1�,SlFH�u!�\��F\��W���&�v^�-�z�1�CYH�,��)����꦳ �|h�NE�h\hm�䚝b�6���d��>s~��D��}�����{�?�e��m=\'��|���8��NP�ǃ��m���b��O�)Qy�:�N����T=?��d���q"N�UG�cUo}$��=ĵ�ۛN��B�������!�s)�M�͆	 �v���"�3���5��<�4�h���
Z�ÏxDDO��f��0�%�?eoD�4^�]0'U��t-!U7�ɋH'B�hܞr�SGDPq8��`�����˄@/�O�������7�S�&���]�9����@�$��ތ4Y*&H�]���g#�X� ;"L̸~�>!�䰮JȘk�V\��D��J�#���"äz ���^�F���u&�e��.Y_�Y݀��vA\q�B�U6�������f�C/3���&@�K���k̈́�l�z5o.7be�e{�5i�M�ѕA�v��{������@m���&��oQzEo��t�esH����"%4I(Z7	Qaʊ���)���Քr��&�d�ߙ�Tj��>|F?3;�s}$*��}�:5���K��������9�D��T큉���m"��
'ii���Cҝ$��",��MK���~��,���<��Iat	>�-Wbq� ����Cu� �m�1Z�n6:s�y�����a��ag|����]S��1����k����i��0�����SQ5ȏ�[j.z4f�[68<vi_-��A%w�?�W� ��9�<�9a���O2I�m��Zη���M.��z?^e~���u����Wэ����>��Vv��t|6����%+7� �상x�礽T$�"���Ԭ�����N��9�o���;�R&�at��MҶ�S���ɬw����	��!HY�߄�(��v_lo
�ex��{M�ɳ��Wp�I�+�$CT��=�"�!�[�_���k���D�*��g��ǂ�Q88)�Gu&1�B>�z����,r<���p��:�vrkQg'��e������;��<������A>�����e��b[�����8uB/�M�/�{�%{�V`6W�c5\����w��.U�fy�C��e"�o� ��
p��(����x�Q���3�ϛ%�!��3�����a����"��<�<���&<U��o��Kj�Cy����8H��w-�/�J��gg�x��j��e�BхH�W�V��B���`NI��J�C�r�[|rC\��]߻�w�r?��M�T�SLuRwG����@Af�U��`Z�`.˘�7c=�D�('��~�p�����-�R.��4�54n�i�%��}��%�K��P��om��p��x	�P�w��K��7ؽ@N�r����!)�k��I�I�궕ϓ{o��g�+1,8o|�7�O��	���d<�hM&WA"��m�O8����Wr=;���-�� �ߐ/��u��{�s=F�r����o�p��*?����m�wF��$�rñ>d��T�tѯ1$@^MK��yL0U��ϙ�}I�	կ���p��KUř��xh���E�S���� Ʌ;E�^"���(�6� Ӧ2�}Y��<��V�<l�Fh�o�u����?���s)	�c�db��K�َ/9N�d7`�O̡claѡ�H��P&��u#,���D*��v��<yܧ��.km_�sI�5��q�VK' ��Glv��'��멬4\{V]MH�ƭk�u�ė+Ӭ�`y�8x���N����9�!>�ZyLk8#���|�B`��f�� ������ǹ�K	@G݇ew�Z��_u����}�\�mB���������cI����3���:F{M�#�`Q�x,�igK}]�P7+^�Y��,3y�@ ��f�
t�ZOߝq�0?銙�r�,�
�bY�V�&��G�|om���r����An�����Wf�$"�h q�=���e�h7��Sf�31����
CK;��=��h��d��KA��������R�b�M/�+���tέ��J����G���#�fo>�_<� !:�1�D�2�� �g�s�~t���[t�4S�W��\\O�d�����'�4:��9�)�,0 ��Y�Zv8,���ҬX5���x���Ǖ���pS����A�be�� �����>�QP��(�	h�fB?!Tء��)����Lw����'��Bk��N�h�5�E��ZN���hڷ_ht���|a㾍l.�7N=��ښ��<wKM�'�6�I��o���l��Y]o����F��p�6�pX{x�:́���u�v�;�s�Ȍ��H�ډ*������.,���PT��</����4j��|�z��l�S�}]q����t��?��������,Z���B9T�W`�������A�.8 ���=���"�1V�
翏Յ3]N�:�Q�ЖF9�k���jxGD`xK`��3��Q�g3nU��ٱ��N�<WmeJJn_�
�n��1�ᮄݺdY
���UO��f��hg�\���ͅ�!�_ű��ňw�����mJ��\���"#����?�X
QD�r� y����s��
���M����Հ�d��Z�ԥ_3��O�;�KZ/��R�!r�t4�A~'�=���Ӣ���>"�0҅\�;����y+�bR�:�8M�'�I���>LO�#p�S�$�7R��)�3�I<�X��?�U�����|�O�� ��3(�=Oy��^��69
8��?�+}�t�q��G'���J"�V�\6N�*0&�G����Y������Z\�&}��:�+��e�8�BF���D��/&C7����6'O rԷ�2���n��.ҥ?FU.G��<O�K�Q�GEbw<s만0X��J�Vt�|_��D��J%��\� v�@�EL�vXlxV65EB    9d82    1bf0~��5�#����@��lhR�z=�9���]?*+(���p�prlb�������v[h����PZ&p����z�z'��v!��uA?��r���=p-S�����u�es��x��}`��R��F��&܏+�{eR�K?����vu������ �pA�.8��y�B�P<��&r�I4���%�8E	~5zN+����a��4b��-��o4�B�����呵���lx,ծ������eK�Tq����� ��O}���'���,�r�'��Z>�83���1������b:BC��n�AK2��"�*`�W^;��Br�wd^5�,���[G�<78`I�-���v��&)��8���'�0�BD-/��ɺʶ[�]dQ�3k��	�5 ������̐$)<���� ڄA�e2�
'�`x\y��R�`���F�E���#�������!o�w�oW�2dV���S��+
���h��76���1�v��
�Um�4I#,[�5>M����C��m�lVx.-C���/2&(�vkbhaW�ӆoJG�i��_�������ǿ�l�EfUO,cn�[�􋤹%e6֥$x����</B��m�.G��O3��Ca��?u�E�@�ă��>���:������0w(�~������h�v�;9w.���s�4�y�8#
��噢k�x
��0��Z����[���!!�]��ñ�g�R>y�n)g#c���0C�p-�~ݣ�P��e�)[{���(� ��x.�CXH��7�-6��A����W�u��_�V�?�Z����YB}zL�rX�Qgȩ�c���Z���};l�7}��V,�$@@�G:�ї$�q���D��|Q2��S�m��[Ӷ��ú�t�V;�B�PNP�X����'�4e��W����� j�*�J��n���j2,M�W�ѷ���
�<#������ݟ���������+�y�/m?���-1��j�~�M�]�y?�sӡn�d�<�*�ϭ�l��c�����3�8��N� �]�YԮf�l>;��@�(�����Ԉ�U�O��}	���)�v���O�e�P�Li�<��c�@.t����Oo!�e`&[mԦ9��3���i��d���t�����}�?���Q�#L|�E�R�K�\�������Q�(Ӝ�z�/"����|�}�?n����7v'I)�I��\��uF�ʸ����g�Q%���! �p��?�ns��� 7s-͡)�d����RP��K4lmb������AX�НA���KXY���R����h��Ʒ��8-6�D�݂�7��#�&�.�g�}����Xۜ4�+�֋ `���	e�G�bE}%	��wa��`\KN|��G�w��
������h]l��aQm�R�}9iU�ꀈi^%��`~����չ�G:B��S�DK�܄��Mh����c���swtO7eU��dl ϟ�y{�J���Ĳ������b?{���8�`8���뛀N�p�Yp}�x\h�+[&�(�헔֩��A� !�xI��Sz	�@�-L�}_U�~\��O�
Wt��=h����Q�+CZ?h9��ʑ(
�21�w�ȘIF����X�vdf��M9�'�C�PI���DRy�t�F<F���=����,]4���F��"*3��C��S�MÆ�509��ͱ ��`�`�#U�F�yΛ)o;��ou��>�:BVt{�Ҝ��"}�Q��"�3J��J���0ʅ
�6��m��O{#�>b)lywBobD�����k���μX42<��PZ���F����8���ЀؚN|����{�����ã@+������0�:������&Ň���hc�[W�E�>z�G�Fpe�� ,	[H��w���%!�(jү/[0��w%r8[�X�h'���ODf�9�l�2д"{�fK�S�4�́�|���o��ok{��?�C�.�3��QX ��j>̂�oj��A�z��k�Y:� �5r��|b@DJ-�sZ��i�< �h������-)��
��mȩ���� ��r��P�v�k'����<8�9���M���r[*������`\�2̥ea�� .T�����2lc>�������B @��-��c��q�ԕK3�z�\�,u�A����.S��J&� ,�H�ٓ�Ǒ�n�Q"��gk���}���	7�q�mz�������%.&��b�`�ce8V�#��&Nw`����f� b ��Ό�@*'�(���l�[>Z��8ś�SA��#;��޳Nދ�1����#UR�������~�R�X��`���Q�b҈�����J�p�����r>G�����܉Ew�
o����HJ�%e���1VGi��U���J����~��`jf<ۗ�zW:/Ƶ[R����sc��J�P�W;L�7s��}���HI���Q������f�)��H
�G[Gk���~Rp�y��[zE�~��3+$>��r���+�6xU

7�I[��3ime�/����<�7�)�x���nn!R���y�@��� ��G��x��}�іy�`���ӣ�No��
rD�^���l�-�]*��j�=�U�#��yt:���Ҍ�Y�?Qd�D3�$�X>-F����P��D3�Z�"=��3$$�˱��8l����C.Zg�H�%d;d��<~3Z�������!�F|�R�:
�t�i^�D��l3��A?In��G���%5�W8����������l��%��c�4*�����KG*��Q���C��h�����g������Ƅ��R=�`�z��1@��o�t�1m�l�nn�*�Y-����"�ٶs�����tX����L�,/��+��|� ��V�9sD� �������H�+�{���9<�c�E�f�ر����2��o�M��[��V-H҃�+�"���_���qlt9�¶˫�CE�Tf�����Ľq�	�<`,���sa@3Aϊ}��t�(f����p�i��iG�
��I�K�l� ��rh�A������6��!ba8X��o���p" ���x�HB-�Pζ=>*)F���K�g�.[� �W��s;�vB��w�6���� �N/����_�T�#�H4��1���3��é�Y�,_�pO��Y�sㅚ��AZ^�5�E|+��}xKI��oLd��F�,�7�X ��fm�i��Ե�f�����`� !c����\�!h�ɺ�|D�(���u��ts}t^2��kI���� ���ÇzTiVʆ��)��2�oƚ�?�A � ���2/�N�[�^��a7��\�&jIW�^�yG�e��ъ��q�i��wqͺ�����oe���OY��zoQI��:k��gj�e`t��&�3Swώ�;�R6�U�2��y��琅6�H�%v�z�oR������յ�W�	2����G$��->)J_s������F����\�L�=���ap1t�J�Oh�R�^�\�Ȥ��E���{ߴH��m��^i%ϣ��S
v�ٗ�u+�f��0-7��w����?�2�^���N>oʊqMw�A��i��B�|��+��@lm�BЋo����R!x.��1��ڙ(lM���x��㿉�K�����:�w���a���\YT���X̠jx��jy�$���ݯ>A~,�\�8g�L?���V�W!�w'�3h������9�
Q��y�ھ�lA�������ͫW)�R��k1�+9�rݜ�ۈ��㯖$ŧx�������.]��О�ĖO���֩4�É�����wy��3�뿖��م{�=�����]$�1~gK;�٥�!OPq� ��M0�������X^�)F7�p,p��t����X�6���u���/y�\+6�㯌��7�H�8��P��ށ[���%��΀�q

X�������⡪��/~b�%H�5p偒��Lk����拿#h�JR:	�L�(�&%���c� 4�rB{ ��F���n{a:��gG���W��c�Dx�0���Q�P&����oc�U�K5�#xjH�?p<Hz��lVUE�B������ܰB�Z�X��N�K�ɲA���^�By���'��׮9 �jz@KNI�Q)|�Zʂ��@��P�����JN\O��������s[��b��	��~�ln����-(�0�/��3z+��5-���#]k��^�R>wh��?��$��^�ռJ) ]�sI�x"����k��'tn�u��W�ʹ2ec�u4@r�+uL�<e�M��"����՟�VK�谂���je�.����N����6
��RBa�bqC���cN�˯�ƙ�[��~[8�甑[�va�U�=\'�����JZ���gɕ%2��>��@�R�d�7��F'R�;�����3M��U|�'�g�ӜF�j�V����R]�i�͗s�|�,�rqm7���R��hiW�(��/�[�<�j""w9�L��Ne���м_�n_[$n����I�v~�HsM�U@c�]:��B�T���������&�n����l�?��ĩ�Z��3�5� �銗^��:{[���}P��jh���Ɓ�JU��-��_��ub�+g�+�t��yW���~_B��)������F���[�ԍk.�IkٷQ���ŖQ}o�:D%=�])�17I�F&j��[�n�t����<mӮ�$F��d��K���I I��g$i�9&�ؗ��iP�>L�0��xջ/����|J�t1�3�tl�YT�Bp����u��o���';)hs}��<�L	(�H)�]�Ճ`��|	�Am0>J��傯�[�D}I����W�݀��r�x������^��h���u�1[�-�\0#��0q��~�,���s�k�yw��N���AjYj���h�(�b�]��Qܗ��H(�zB�d`�ō��n4R�kLa�Y"��Փ�<R�/����
���A�;����X�պ�G�c�O\�푍�?�M\T7^�o'�5�J��Z)�e�ې��БYb����+M�J����>�q�'Ї�_gR�:P�s�7��2O�T�5�
6�`&����2C���!w֎W�6t9ըT��1c��xJ��O8 6�X}�����-�&�g���+�����Z@��/xL��3J6��=�毫]zM�+�_ptt�'>q��2\@�����W	2������a�6�=	�f�
�h�'�v5:��&J�~��wD]ṣ�hN�]����Y����ЦZ�7>��!�Ɂ�yX� oe�=Zdq�:˽��k�&u�:�6o d8�v�ãsB��r�V��Vb(ң~�L�?��ԋ7����s�P��uI��3�s�}
�u:K�	g���m�Z(jK>z��7�i!Z���|�j���W�a��Mf(���ЁT��g��#�菚W%!v�Q�%^?������ۍ�u>�Ԍ���CKEN">���xw^w�=CN?X4� �垔��<�J�e��Ɋz==2��r*/Y\01w#����](�mf��{x5�ҫ�_ү}��Ɋ����gA���P�5
�.�\'7گ�P�S�s�^�4
�^6�T<���fN��8�3�q:��_<�J(�j���U突������Na_�1!z(�����m�U}�|�V�X�s�sF�)��PRo}�ݬ�p;�v�Y�Fp���D8k[�:��i����j(4�������
9���:<��q��gv�����Z	'F�].�a'1��%�zܶ;֋4	n[���L��đ��G���9)c���ChH���Y�]S[:oL�9*��K���;]0�������[���p�;gL�~Ha�e0S,�sѮ<s|�~��p>Yo��}F㸚�d�e�٥o�2���*�d�	�C�9��	�޽k���O�Sȑ3��I�ᐫ���BS�U�c����|��w�N�JE�v%�#BziMθk؎&����������fk*���i�Ƚ�/�W�0�/���
ޗjV✱W�њ��J�k�B�ZO>�`U�}S��#�O��  VPu�B��JU�o�=@��Y�T�N<@	�V2\�iBO�z�K�ɼsȠ����hH�����X{�DGo����1���t����	Mn��& ��~�}J�جBI.��} :Cbbh}"��;�И}�:�����i��eq���pr-m5}f!�����I\�|�����vQ�~W�_�͋����r&��0�!����XOK`n�t��$��zJ�(��*��i�鴊I�ܐ�E�+mR�@�J�p�����+���@�v�ƣ�x.��¤���'�^�ՋH���v�*�+q��*l[ת��B������ ��B�^|}�IM�"�Uw�[�"�*\���3Ys	�P?�5���' �4�I��p55��\T<-�g	�m�%�	�Ab�>��`�TҀ����Q�O�� QU�=An��$4��B0MN��K�S����Η�h��+Y�.$B	����4n�����$J4��98l���	Zvs��K'2F�ue|���B�FSxP@�v�~���[�z��T��������/�͑R��fVOW)��K��@�f�%YBs��ٹ;�$�E�EH�MQ��	B�D�N򒇏��2+6�՘��ˆ�qI�ܞ�^���G���2Qs��Rv�24h��2�H�;����l��A
���|��oEL��+U_��n�>0&8�ڶ�e�h�����Ƀ�A�  �j6���ݳ��=h�5��;1��K�H, ,�4|�����Mc��M�E'��O@�4�(닏��$���'q�N�oAX5���%l��Ph��� �f��ԏ��ڣ�J��dB�?��G3v�֭�3��j�z�_���~�����*�0xP���:f̝����&⡪^뼇.����aǥ-_��`��ͪ�����B.bx����c"@r�4��i�����n�Vi k�H��*�����J#0Ȟ�}n�D_ =c��v�폧~C�6�E�A3���Ԉ��Q�s���1����D�2�-XMqu$�M�5�g�9��C x���Ҹ����׶k=��0o3��E��nĮ?@4=�g ԞݛT��;�W����Bh��Ѵ/_c:�j�t�(���˹Rb�:ՙHX�|
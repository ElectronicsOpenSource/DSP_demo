XlxV65EB    fa00    33a0� ��ir��g��<�����Nx6
ք1���2��kܴ�Ci��~�!���K&���\ʩ�w�kC˨����پA���yZ����l�v�b����,v�q��z���݃+�1l:�n#�P�:O�	W�ɚ�SB���DΉ��7� l��8
�EZ����_�������Gt�h�wƹ@/*�����X�i���x�J�ї�!���&�Tg��W�7��S ��噎���e���c&Y�F��&�᧻7�@7�ģF͆�U�r�M���"�C2P�M��I�E��.ã��CR��|<E���>8����izT�3����wG�cn�Z���O�K4�%Ɏ�T��A����S�^�3e�I�j������ы���s��AE�S�3��4�� ��,��@	���a*I ��/���[;2\�x��� 3�� \�H��i�#F�N�$�M��7T�G�}]?o��sk���5�J��]��\�'?�Z��Z���&(l�zK˼J�2�&C��*G.kŮ��ϊU�������Qg��{<#��W-���ni�y���@Mc<�z��`E�J@�1=a0q�,{YK,�֠=����o�U�ߢ@"��Ο~�HnJ�]�º!��o�<:�汾NT�/��7���Z��!:)YN�� G��Ŀ<�]��+���`3F�p���:���7��ZO%x��0�5ř��|��\]
��
�'%�u����"���I�<06��	�s�5����wV4�K+��)l�ϗ�h�pOϣ}�����A�u�( ].I�7*B?/�������:��%9�)"P�m�����n]kM.5�`�ET�̑��sɚֻ�{��I�K�G��Q�o�k��߰���O�97�eX��U�R:�L�M<�߁�gb����c}���T�>�����E�9�l��������W�=988s!�zp3�Bde��|�	�4Q2���ʂN$��%T�&�լ4�I���p`�$G�"����]����G"�������Z)�CNӁgw�E�����<�� ފ�ߍ+��{���m���D����!#l��E�ѣy�(��z��3=]	�lV*O?�ߞ���H�kg_�څp�S;ʼ���O��!`A�-�EƋ�鈑�%p���z/�v�W(1��e���:n���x�$.��[T`�btH�~��1�w��`&;2$�/� <��S�s3=�I�_d1��
�>D�0�Nn~5�VA�D��TV�T����^��w��Q�V��˰PH��p#G��"������g��aH6��|dyD��b�e�$��g�aL��g���L�8��T�Eg��YE�^J{��,��$���X}l�9`�O4��L���?�m+�k�mi�Y(WF��K,�? ���0j�6_�5D��^�����_)�U8��	N���%�SAO��H*4yO>*� '����v(y&�7�C��U���kΩZ|���9�3� k���f�m=�h*�ޢ0���+����WR�#��� �W��{��S��^@�d����{-�D����D���!4ul(�@FTi�.��	��{��;%B�����>aYX>������]��i��a�D��KXƁ4�\�Hd�I?���E��uR��-.j�u��`Y�3�
irU��mN>�������Q�p����ڕv1医X�:Ya]�2b.�����q]�^1��؁��9
u� �uU�A�~��٩�
�
|�0�{�����i��և���U��n���X �����H���ƖqJeq.��Sg�����Jpb?�{`Ff���b��0�k�{��a�f�M3��M�0l�b<��~h"@��R���u�f<T/����T2*F�����&k4D)����N+����߷��Q�8���K��Y�7@��nl��&����W���$��=Ag��p4H���3,�O;I���M�R�Je\��WU��4q�����sP�E��|�$B������C��؎?����Y
���X�=�7��;ՙex]H��̘L1(� �\��­��|�gR�[A��_�=�\�h�'�5um�zh�_A��ܘ����������R�a&F��� �l�V��U�W��a/����� �l�	UPG)#���m/�����pZ ؇	��MMW�&Z��Ё5ń�S�V�`�܀���4��F��h{H���I�r�����P��a`o4��1��� ���;��N��p�ju�[�-}r��2Il��ߊ���Ʋ_��^R'�8�<�։���\��T���	��ޮ�rZ�Զ�I�mDr�&OQ�׶9��5�߻���v����+� ���ݮk`����i��^�.c����K&�""�۴��T�e���=i�8%J'+,"-'zĂ�:�/IX�%��lE��;s�
A�o9r}���¼�ƚZ�Я������J<���{��V��N��d�[NreU�C��l ��e����+��=B4r�l�T�k<?��7>@%�3v�q�}Ձ۽F�=�jA�iz�]�7��8�A
4����ǰCĖI$4�x��-x"���s��Vq�5�AʆbŌ���ΰ��d���)�"$#�UQJ���4I<�%f�V�Ox���p�QdpQ�����Z[Ŏ����|�~�RT����0�)u�ւp56bk�Z"�clȨm�:`c��LP`���b
��1-n�,�ɓ�aO�2~�� ʍ��ɪ"��YI7̅��,�{?�.�y]Kt-֗�yn_UI�䥂��	+�&�ې%mA�1��"�@�~J��np��	�¯Ӌ�m���,�?=������>h��UM��rね*NZ ��D� �1F�Zu�y�K#��61���dqI�KJ$�Rup8JZ�ІΙ��%�0���+�p��s}�xc�ARW�$인j�UV5�ܘ���wc�s^�h���j�lz�m��z>���I�`a�ɖ&�uT�}�
���B���0`�������JZ��8|�����c�̛��R����.�0w��-�DM��Y�`�J+Ke�i �D���_��X�m��EL�?ŉ��)we�s�A\Ψ�'3}�}]��Q���q�-v����e�<�+ a�f����il�h�C�=�Gk��h9��x�
#5 �������c���w�~~R�qKTE'�{���S�N��u�V�z!`�H� d6+�o�7���!�H�J�}^��:��
�����σ���y�#�TE���~�}���ȟ�����KxVd-b�����,P�k�𘢥����6��Aq`_-��E��/�鏱�s�&�J�W.S���A���3�T:�'�j��f�7���|���3Q}��-�!�t��gj�-Q�zc����\�A]T�ݺ!���TP���g� ��F����W@�&N"N���-Nw�zf �9.h������|K�8��}����u��xZFoɯH�ؿ%ӭ%�1Dqg�k=������_8��[��7_i�d�I���*���
�[�e�Vo##�ě	�c�,R��w��^v���ɲ%�ovF����/ľ�Ǒ��qɚN�3<2
��ᑙ����\%׳��e�_T9ϰ�&�u��͢P����o�l19:���ʰT��ި :�In��V��O-���`ہ���H�����K"ȷZ�B*]�HQ¼�����L�q�cFv�-ş˓t�`�)8����6�<Q�m�0�8F�d��l�5�,�L+�%��@�M?�:SE"���I�W�G���3z��	J�@�Ck]�2:�Ѐ��.gyYG�W�R�\�����������%�@��mɟ�LH鼶|�M�]-�r�T/�Yr��g7^�����dC������L�ڜ�i�c�/�F�t�Lsw<{Ά[�p�(M�h�f!L�(����������ǁ�sտ��i�$J�Z=�_��Pe�K	��l�u�+z*��lx\!�����!;"�y���ԭ�d��@�Ф�U�y�Y�!v��Y�)_�c&���r��{��ީP��|j?wMRډ����aJ�T�Z�wZrI��XD�d����u�C�x؈9��j��� �-b��;3WA�5�v7���*9�زj��G���@���{gr�&��c���L,�� �����S<��S�e�	ч[$���^^�A:"R���4*IZU ��Ј���H�"%���Y	ܯ�5�}�Mp����(�	T�CV�+�r����0����j�s�����C`l"�#0j�d1�
�n��=��	����c7�}��0';��#��P�=6����)�=�}g5�j�1�w��LöA�̏2�ݭ���=��^Nm��Br�`+����:���]:#mY��#Sǐ��(B_�O�J�5`S���]�9j�Rv����}w�`	 %��c��0G��G�;d��Z_�q{@0��OuV�u�wW���l���p��$�RR�4��~� �"�k�!��.!�4�n;��Hؿ����mk�l�� ��d!>�ͬī޹�ڵh�GE�>�s<��u�L+w�Z����|9�[��Q����cf������ �Rl����O���S�;����F�`��Z�ԼN��A�Ij�񆔇��Z� ��6v�݋�����&���Nv&;��8�<�`42ݒ��LE@��Aܹy�pizG��O�YѳuɎ#�a6�.�o�y���|�؀��������tE�0Np���h���E��n8b��5���
�K������R��Y��*�ZI�D������^�+8��������g���2���?rZ�o�_u26Nj���8�;}�:6�ʟ�נ�^�6447$A�V�:�p��[�,�!��(5*�}��7r};.��E�M*m�x���!�������M4v�+H� [Ďd��$[ɏ�?�FI�3>]��*=����Ur/#�ex��7��/ ~���ijB��{ ާ�s�i�֧#"7ܞ�F���կ���]����F�^c�$|����,�o�ǧr�!�+�c�U>��W���P�L�n�Õ�A�;D�U�/�H�k{�_qy��z'�&W�g|�����<�9�����.���+�q�Sܥ��ӵ~�޻�U���BD�ˉ�4�^�g�=��3P��<�2�
�n��v~��_{���{�4q�,ց_�Ą̎zh�Kq�e�u�=kn2�r����gqq@8�J��_]�/5o�TSs��3��&"E����h���pw�a���L�� i�v����A��پ�������u�����;*�|��`���=Z*�I�wo�[//�-��^��4v�!`N��PyŦ�i��,�o�8��<��w/�g���z�Nz�
�����v��h9l�['B5�}�/�M�u�i_�v��ߎf�m����f���uNo�sV�J<���+ε��Ö��S1�'��ᘖ��&4n��GSJE��P�:�^��u��ꆷ}��3
a�X.��Kǰkbt:eG�*V�������*,��n���+<*�Y[��$0����ݟ�YY{�hŚ�@���dfkv�AۧH���P���N�dxt.ηQX��Z]`�cP��h���U��^e]��m�0(����ܚP5��{vY޽{�ţ�K>��9��N0`��]�D�(C�����\�ss�t�1��)SC�9���0 �G��ט�ޕ�Vw&��L�b���z���z<R������Za����bt���$��{ЯJK�Ƚ���5D�5���oy�	]3uϰ�D>#�D���E�V�� ��V�D{m��CD��Wͣ����'zϑt%u2�./S
���n7�uOå�3��zX	j_@f�Ы��Oc�'[g�Z��ߓ?�$x�����vҳ� 0�6��>�mQd���#��q��i�U���*�P8��1}�jI%�2�}k��U�6�ubr�B�x�T55��2��J��j9�Mv8���b�K`��!M8���}�})հN��-ñ{1���w-;V�����I��AfD�$"�f��i:���g�j;�2���h����!/��=F��i���F�:O؄i5�W��&����5�����tm:��\�5��<T���l�R^�i*��Z�h��JԎ�E��U��m#���d˼�e��mF"�����Z1d�pǗ�������!A��9k�d�ZR���ir@KG��@��-8�w�\`�T�����Q:dV���bd�8n9M�q�9��JL��*v����(T�]=z�byRTi�Ł�"��βl�.�Z��e,ޝ�)j��?��eXg�B��~����MUp�pMPWf/#�Ű�e�!��f�1��� �a��mU��R��O�gQ%�m��c-��m�C_��A��J�Z }�5�*��~�'ν��@���o������G�-�e�OC��mC��b<G^`�V܃���7N�L��mÅ;����F&PcO^�'n��?��������ئ�R�ʑ~��"�f�5|���`Jl��y��I%�u7�a�a���`���]�.+�:a�+�~���4@)�G[HT�qM�)]�i�79��qT����h��^���_��gX����V�K�4GT��>KI�ea�Zi�3O�k �;�zO�j����֙b�׃���V2� �)�2�gY'6������cO_�|�1�?�夬�.��8o��Q���\�b)6�}RS�iǕ5;�:����m�1��ԃ��� ���G���|y ;����W�t����Ɇ'C�Z#��;%��X����E}��G�/�4��Mc�R �}�Z�`X�ؾ�v��� g̬F�����2�1��b����\����Za̚4x��?������W Ϧͻ���z�̯T�,�r������z�����/���#�a��.{L?�Ѷ�h5�Y�Vc�S8��bO�S��~�^iԸ���؍�x��5��l�Q������.�1��J_a:,�`$jÜ�x�~idc" �H2zM �?��=!$���N������W� ���E-G�����[UP ����M�=���$��+���=>��ip�W��$̥��ֱcr`.���t�qO�?8pſے�oM�`�Y8�g�����J�n�VH7�"v��.%�D�گ�s����[��)!�wD��v~+w*�Ѯ���(���)�˜��X���7��Y�D����s���RX�?�j�����S�4\m4��o�gR停ҕO9�.���Vݠ� ��wRa�TF��Eg��@�\�p6�tGƀzz,�4��P��(�*Ą݋�����<�%Ob@�����˵�W"Z��i��o�B�;�Bܕlɸ�{q��̰b�3V�O�UQo@L)H�L�ؤk��"�8��Q��~�Mn�5��B�U/���c��%���]Ù�}���v$s8�nBZs&f
b�)�wo\-bd�D����ӏ�[5��֝�yY�x��{�>�V�|(W��q��4����}�ͳ���a��J���7{$0�9 ��'i��)0�!KT��a�!�"�%+�c�L���{��t�wK��Rl�.션K�?�=I����K���]�̜�RcT�����p'���J�5�AP�R��c?�y���^��Z��76uО__HZ�B"���;�1�U|c�|���,t��L����c�I.M�1��.m+R���2'�ȕV�)t'zs3�B���hh�����=��[�O���H����+�}H��ɅG��)�o����~���t?���T��:P��bk�4�,E�)�tOҮP�R0mFέ��S�O�Zv�?M4�Q^"'���ߥ9s���_���h��{n��Ռ^�xl�P�>¦7�'��c�I��l������h�é����5\�yڦ-ӷ��*�g���RW*l[��(j��+�{���2���[>}Z~�A0� S��:�K�H�T�٢�["]��>��?�/�hS��xx3��ۚ5�+^>K�����ɟ����ߜ:�L<�јo�t��Y��q�7�?�
�s���c��w���N���|���\��H����s8$�]w,2�����q�A�2F����O}`NM�N�߁���WG	���"|Udw��:p�g�;P ��ů�+������Ms)|_����@���k��L�*g�B��4�u
����*cR>�M���ꭉH�WV��Ba 1/���g�p�orn�U�q%d!:��N.��щQ��_�kiCL�)Wb�=�b["= �GBɳ@bH��JD��=7N�,�Z����N����0�C��m,?.o�̷�b�/��O��L�������Ά��#�ds���#Sg:*�PmI��gĐ�@k1|8��("&&A��oh�=�u�n��aϜ�Y�b�G�N-=�Sa�����L��M��CS,�X-F"�Bn0�/G�@e�O|���2pyy|�rskb+?a2$�D	<p�*6h^-�T0����'&�;Iu�S{w@쮌�����i����(��k<m�(��&M�Ei�)08�`>{DP� x������)�}��@��<��Ǌ��JF
�n2���ԅ֊'c���N��a0��,�Ÿ\�'��z;�HX���p+���ڞ] `�b7�l��QE���=o�du�;<��2�XR��w^�2���U��B�z�	bo8�0���h�T�ۉ���Z0���t�[�1ĸ�����7��$�������K�h� ^+0G���2c'��[�����ާ��!G�~ZC	��P��M���{��^�ۋ'�G� �w�f�wp�_�ᩤ�>w1��ö��'OɤF��"����D�x�o����o ���5�˒��;F���0�������A�������׆��m�t�l��OV+��#]��2��6�M=�z�W���E^���6= %��2�t���<�Jĥ~z^�U�y�ƙj�2:�f�"�Z.1~��唧���	�mjɬ��?ΜMDDtfw�W;/��d�X^t���'1k&��
˦k>��'vs_����Wr�R\���t���\�@)������ў�1��N�4Ϋ���v��נ�}[�e3(txc�dG���ֵH�J �^.�g&�����Q�}����KV�|�v�����t�n�=�e�s��	��Dq��b��A��5|�$]�ǳ����%4g��J�>8ec]�`A�G�Ƨ��P����f僛�hk�5<�k��z~=��j��C��^��f�{�k�d��[�dP�[�GV����Q��f/� ���xѯ�>@Q;��^j��(���o7�-�t.������8{j�1��U�;�=�t��EbM!��]X�Cy�u��o�9��a�j��W�$/U+O����N+���K��t2��#z��A�/?�<d�����\�Lm^G�^��Z�����I�[�u�s�B`4��.,���� m�6�PKq#�(B!��;�Oa�^Y8g�w�xK�0�4d��)r�IL߁O��.ǈ���0�B�|g1w�x��M2z�<��I!�v�jrdf;wL��S�i�����q9{3X���3m��_��S����DNF��Vvj�����Üm<&<W�l{�.�m�0�oY�$d�Ҵ�����3[M�I�؍�-��s����&����|r��jCt�'�gB��]��Z��rM��.ҋ����7�ݑ91��^�����zWh��ǑC�z��w�\�����U�ǝZ�+Y-��!��/ӿ�q��	���db��K�T$&;mh�ߟ#�| ����y`��B�z���?��%�%"U�"3��\��,�)W�ꋼ��)�=.��?���'P�͆`����B�Ơ���{�|�k��Bbck'ʻ��� Z�p��^׮����&��ܻy��y��d��uӪr˖S7<·vלR��aj�hP*0Ƀ`�Ta-���;����Ecͤ�����7J�C�g�QS�d�jg!�P-���Sm��� "��OEce����[{:3�.�
'��h`������ñ�N�­!���9�Ǿㇳ
o��?����޶2�A�kQޒ]UJVm�'9�2�Wa�
�>�/���汪�|����s>o�"|�$�ܦ��=����e�벳�rk0��u+���0���s��.Ovm��-�>�h��f�ֽٟ@���(�B���jS{&�jä�)�,͏�mK�:7����K[X|Y��~�D�[��� u�sh[7+S ��
@]�:�ZF���9����?I��b�������޹�z �\>%����?�����'Rp�{ߖ�*`'0�`+ő��pI&*�	��-U�-r֝&�ln_d�'`�y���5<;]�/ԕ��%	��|����x�W�����Вg3\��+���ʴ�	Ŷ�n�ܱd�EE�5�P&�>~�d���JJ��(�B}�b��_���5*�����w�SB��3]ˆ�G@m�}��{g��K����t{U3
OQ�1,mu����V8����L��`S�����>eFQc��+����pπ#�Xv����L&^б�{�^2�aqq����z�ע�q/���k�e3�%��x��*Űf�!�Y��.֯���p%kv��}~钴��e	���,����^�o����B1`|gx
�LO����m;�*<t���j���+`�I�\>���p�i)3�HE,4TF�/��Znr�v�$Lު��/�頺��M����K�U�)T���a�D�o+9��yA�;�*S%��K�ϗ{�W�b9ٔ�A%#�Df���EXqw\p5I�4�ޕ��W1�j��9��q���2��͡��m���z��f�E�>��p�Vs8t,�yN�lh��hI��f��g9���h�[Y��C ��AD!����A��X˲�j�c�.�\��X�wY��7�~D�{��1a�iA�n��h�V�&}��l�1�G����책�\Vд<%$��q���� ={E�$&�a���&Y��ݾ��t����W,8������8��zG��)zj�2�����װ!��&��P}���YY������8Omg%a�i��|9���*�2�7����;�~��T��a���+%�y�,>�r��06l[NY B^Z�kS� �WH��iꟑ$<Gy��ޮ�����hI��#<��� `]�y�69�C�!	��<�ޔ?���cNq:C������9�>��-{Dm����j�2@�7/X��</!��k8��a��kG��Dl�4��V� �Q��>����W���t��-��q�)��Aփ8O�wȬ��ͥ��; �l�>V��`�b ����%��Y�%������x{�P�$�!��%l;.eN��Y"�8��٩���a�C�+��� R�\gB�g��:'k�����}@T�w*�&lO��A'�� \���T6Š�ut��`��&�">_r�A�ۑ�O��G"��A�B���G�蒴YT˕�j��!:!�y��������7O>�|��-�0�����
���㆑�E�D�G��ic�>'���8����?���x}�<]��)y]Wr�r1� Pκ�Y�S�dk��TʳJ�w�8��Z�tpZ��/��\Dz��%:�i��''h�陒=k�`���{���2�%|'i/T���xx8�?	�6�M�����m�.�'D�w^k
FՂ�ۚ��^�ܡ��"Y���0��Z�qxJ��-�v�M���t{��އ0���I���$�r�&ݝ����?$fA�aeԳ�}���L����C���g)�#f���ء4�~0�yPܑ��@�bF�L��W(�I�4�nyK%J�&B��L�n[:�:��nʻ��)F����^�Z�X�Bޭְm�At��PI�6u���;�[B7D�6����T휝���Z�K��@J��c�i�&6�X�\up+�%�·X���J<	��Q�&���_ɉ�so$������`sW����(/��.��I?=��g��W��
��|4|ꦉR�>^�6�$h�}����A��n�N&ǔqU��� ^`l��6����,����*����f���0���o�w�$+��2�9�/�d.��So�
K�=���AC�G��Er�y@�հ@��4�����7w�4$���t�KH6�K����FdH�g1��������A����+���$�5��q5����HD�{{�
E�{L��U�ɐfh�c��(@N������Ée0�o��x���=�a7AP~!���H!u}�}��]DU�������r��Am��Q�1mSs-��gGi�fl�������@��A�����NS�Q���rA?Jn%6���˓"��)���f@�^� �qb�p���8��j�;w��>�w��T�Նŀ��zw�.%
�ms���j��7��؛}�>+9&�"�����.����x~I�wJ�:Fw��J��g~r�8�g�{rI�ݿV��k	ۂNb�����ڨ��}j�#������r0ݔx	1��99q^E̚�y&��pj�4׾j�;�� KE�K����"��!�u�'A�_q�d�X*�x�3�yg4�0":x�~�]����ןǦ��ix0[�z���;������O�V[�M-ay~q_?�=I�*q��*ON�q��&�Qo����8��̷GA���=�ϊ1����x&,Z��Wx���N��ya���sC��ªo�]YV��(���}�A{ B?q�ݟ���%+����rGU����\O)�N����b/W �)��U.g�#Mh�枏!��>7$7�qE]�-}[<-=^L�}�61�ԉm��%e3��ɺv������Ҍ��e�P��|�y)�
k��Wf��[�?5[܅���h}F�3�y�;��6��%o�e^�B
��(���}���Y�XV�'N}##a׈�f_��EFS@x|<��" {���sLbpT�}���BkĪM�8Σ!�h�T��4A�o(�ˊ8^	��3�~#��h�~�~���z8�j8�YQe38	�ڦ��O��N�L]��"Yuj�����dɖ���.�-�C%0/��X�Ø�.�/�u�A��E[0�xQ�
eXlxV65EB    f8fd    2c50��ߕ�6��}/j����	�]��:����:� �g�#i�.A��pq�ݔ�P�H�2�5�#0���s�oF�X�?h�)�,������oo�v���D�GĐRd�{<"X!���!�W��#և�
��}�BO�ʙ?R�~���i�m�� (@�p�Rbx�����.��������s�M������a��GV�!��R�[;_�Km�v�	����b�J���nRK�Ll�}v�ՇOR�����|��� :��{����y�,�U^Ch5�2��q�kQ��ѡ �/�H��R��W{��@�A���QRog[��sAlg�S���;O�H�}�
{���_|�+�-k�A�����\B��8x�!!�4�ר�CXaz�3P�R$�K�%/���o���|eB���+H:�{3NM�a@#�?VV�$ر_l�Z�gy��\�����嶏f��-^ �j���zˇw"W~�IrÇ7�u=�	��N/��:q(�|M��SDoM,"�������J��ЭbT9�sBm�/$�(_u[gf<��)��h�ծEc�-��9���E��V��1��#�tLʥ��J�� ��"�*��k���eۿ�K�����ʬ`�=�D	l,U�I�2�l_�kI�x!��vG�K�};�������0f#U�ANKhDMp�����z�����Oi��ijV܄A�����o+6N*�x���@�.�T�/b/�,d
����r��xZi��l��߿3΃�<��Q�ڞ���R�w�!h�ߍ<��)I1�s�]���bA��M�%BS�Ł�Kg��zz�G���[v�7�J;��j6`�V�;�����z+ ͜�$��P䶋Xn�|b̃Wx}/���73�1f�̀R�MG(%	�,��]8ӖVuk��w� ���x�1q>������5A���ET����$~��^���I�1��:��e)�'KDXE��P�)�HYN�����Mg�t-�� Q�(Od̢6�A���`�*���4�Eo������+X���� ~X��3�Æ��߾^�BGRh�⢯*v8	D��A�ܜ�o���3�\�Z����h  H�V�&aY�4Ҵ��K����r��Ӗ��N!���C��Z�x]s̹ZJ��)�[�1C�+�
[Z�fd�Z�g��tj�#�J����$�H��S|��������аcH؋�~0=�h�XW*�`B�t	R㕗����	�s��8� �H) �%/���re����XA��3���Y������z�z-���N,���|��J��
�O�Q��<e�����$���6�ǰ
~���*%-����,�%���p|T�+;�e��sY]���KjWm�\-\XQ��W0�n�������cM�&A@ �o�[TFT��AH���p;���`��Z��0��,�@P)��������j]IY9�sQ�0�9��d�|���@�^#���B�8��ɭ������i�Z��=��"�G��+�.�Z��r9c@�Փ�y|�-��xŴꎇg�G�u���*D�Z,�&�/��DR��U(��gv*�,��+mi��B}� ��ޔ�5
�;��}�RXY\��r����uW�`Mй2��غ�=�$���5�E�ƌ��p�(rC�+� �ei'&��;b�yl� Vt�����;}ц?Km
��n�+��3�U�T����;S�&����|#����%��K�,�-�qj+oH^0h�Wm7��{RQஐ�l_hv��9)�%�F�9&�γ8m�9Zp��I����l�Y-�ꇟF���n��g}��U�H}ZCY�~Ǟ����c��i�;�_�B�o�?����:���GY⬯ ���,~�5�wh�0# �� ����"k�%s�]b�Q�.�"��~�P�������E�B˙s���1	��i�o�D�K��X<�l:��X�@&�%��>E����[J-!�����/��� &@[U�yЄ��o���vq�{�X�0��0�,���Cn� s�a� x Խ)��^�l=�LL7�P<��(�8�V�k�t�����Pi����yj�;��}�@�<	��*̏��qj��!��y��ퟣ�k��@��n��D^&J�m$���̭�<��pt���sdK���,���ε!ۿ�9~���Պq�M֡'K��Ǆ�_-�n靱u/�
Y��yri��#+Ve�,�z���IRB#����f��9/���U-��b��R��(�+��������Z�P%(�$"3�2xK�?������vX�2�mF�8����Y�M�w�z)P��=��i���pb��e�C;ޮ`<���]�"OLH��Qq��9Az��⇆�������>
���k;d+B��50�q���-[�3r�qMPy�A)?՛�EI��R��,��v	��a��|8L����$68	Y�w���lក���jc1;��	��S��ź���b ���= ��&��<X�P����/���q@�A�`��C^2���F05�z�'���w�����7
H�\���4�E��po�������W���Y�����NS��e��^�f7�|l���A�=lG����>��N
�h(�m�Mb�x�M��C*����x�u4���J�|w��vgߓ�$�U�3�K�t�p�,`$1 -��qU:��c_�⨝6ח�4��Lm6�e�.$����p+�c��L�ͺ�3������e�Z�E��E�����G]�7c]V'VzXU��=`�O��2�����`��W0ei��I��j󆾲 {�e{rv)DF]��F���𛋭Ӂ2ݽb ��rl8g4�j��a>Q��*GB�ف�.H��ۉh��2�i�(�]'o� pӈ9��ߒ�S��8����u|O�I�t��4J4��0i��m��p����5u|�˟_�����B z�l��F��/����PJ{�,L5R�w�g��	�ޔ9D��r�x�|"�ߝ�|x�C)��>�W��^%&W%]��FN,ãz���IH�Ư���� ���}�C�}[}4�UT��	CD�7�`��#��f�Cv}��5�U�h�#�樼�;X��u�Yz�y��@�:6-nޫ�w�	Q����qzmy0d1��
`k�����օ#5:����%���B�爌"�b!+�H�+X�"�
o�e���T
��/����3���Z�����������RY��J�z՞g�w|᪢ς�I`s�i^>�4a��[��J��?0�!"�Ux�3��bb醅���h]���k�2�?���o�&�l���%s�A��Π��4�V��Nߐ;wf<�Ư-h
{�g�ف^�@��e#�$��F�Ueb�&�;�k�Ӓ��G�9���)�A�!U/ꦎ��2Ǡ��nRe4������S�#i��I�r}��,�u4�y攐I�8^�
@I�F�Y�֦�0���*Q@V}�H���/u���7�߄���N�-�B��k��r��+p>BNօW��>7�J��}�ICl�3 IC�M��0Bw���n��ht���Fs�z���^":َ@0�	jȬ�����D����J$�ӈO����!@��ۮD�r!��Ov9��f��N�,�$�E�J�?�dK��`4�� cn����1����j��ex td��}�zN$ɡF��-<�o����9�!X��PG�@m'$�S-���p�&ljlxu��.�[�Ǆ��aF6.�
��ލ��P�N|���R�]֋G[�n� �C���*Q���܂�)4u�K_�ǩ�q9�_�Rbڏ�`�B��fM�90]�x=
c ����*GJM ���o��n�	�e$��|��A�l�e�^�i��LM���ZM�?�����/��Gkc�ZI]������2�{\s�P������AsS�^������I�s�82s�;���i�/5����/q�}��҄�q��'_�{����	��0=G,_��C8����K�В�kx���v]�j#�ɂ���w|�(�A�^<�n֋�`@��_�I�qg�G��x(�%�V���;LD�������m�1۪�eQ�Ϻo�"�MLc�*�� ��d��I=��/��TN J�Y�$�I^�t#<��&F�EΞ��jR����ȖB�'1Z�ղaNL0���|1�m҇��[�9�ݽ��R�i�]Ir���O�'�<�H��S�r�'����&��H� -�;�
�`��[/��������х7���J�0*miZ��<��y*�ҥ���� �g�I�����}#���@X/�ٸ��j-�+i;�M��[��2?p����#h�
f euS�в��7^^x�8�ۯ0��]6�C���r`*��S�ܢ7��U�l��Czrhd����s�9m���Yʘy�J1���P���c�h�
��[�x�b�^���z
)�.���|� ;N.&��I���ۀ�u5�cz��D�?lrt��x��_G��8�u�:��V�NY���fL[T©E�$��]�oL.l�bs������%y9�t�f�_Gs!�D�,,P�q��J�bc�X��vL�/+K�Ju��j_&�Q(�n��aXP~)f��m4T���2;F66��olJC�����)Ҝ����`�6;@��[�j��Mե-��{�vڇ'b]�!�p�����W�>]����6 �A�s�2���L�o�o�=Pel��õ=ׯM�?.Ъ79��"!����r��PnN��!��IB����Io,v��u�����+��'����U�~��}c�����{KS�`t��
��̥��R�(*�x&��<�2���Uq�(wML*4g_��b4�<A�-V΀C/R\B�UD���U��k�A���c�6�N{1��֩}��?aU�x���û�>=/��!��C�� @C�4����٧�de,��I�'�,ldX2yif/մV�dS"��
O�ZN=���2kd$k�J�>'��ot�B�t��F(#�?5N�Ү[l'��۶�b�)��"���apn�q��^�>���2	���zF F8�s���1U�@L� �K�/�X��yX�+�,3kЉ��	bv繱�c� �>>�g%��/�{�/���)+�t�m�6�n'z?���LS�� F�x���Q��L��F�1����i��n"0Js+أq�y�R�2�X���VX�=\7x~�ŝ8`�݄�*̐�����%G�U]�Z:���h ��
c��f�)�pqp78;ۀ�������_�o�����i0�H���2���_��И6�&�5���]n�
��;�9l���]Aԙ �Y!���3�|j	ui��o�2���Ы�UU����?�V&�S~7'�+{w >���1 S:Qg����+�T���(�~���mWrqԱ�K�\|-G�8]>�B�)��]��l}@7���3�U�2����Б{ܚ%��İ�NayϘ�^}ll<�r�hȜ?��ہFZ��5L���q!�E�I"�j5��
K�W�p��c�Р b�*��џ����N�R��э�Y봗i���R�����~����J1�F��av���%섃���\�_�� 3\�5���A�E���w�ܻ+��P90E�C5[�	g�$lڏ5ܦ�p���:�R�lJާ���N�E�_�Xt��{�j��<8�E��2|�������Q��7)Nĵ��8�E`��ڋ�s���T�刘�+�UN���u���í�-ms�_�W[@~�!7ܥ�T��l�mb���?�%�x$�Yx�1�(tE&���6���=Û���q!��ɇ�-��I�Cؽ���H����~�E`b���_�L>��̧�I)do��?B���M���#���ԃ*��3Ge!%����T�F|�w-���HhE��q��dHU�,�h2"(��O�Ap���`[m��OG�_�W�����v��7h�����08�S½w�g��7��� ̜Kq�9-��4�~��
%�\ܚ�M�p<��q�4G&�9(1����#L�5�������oG2"�¢����t����Ώ��w�0����CV��S,�ېa�3��9tQ�qSHqV�_/u[����7�1s�0Ж4��Ѡ	[;�3f�L�lrl+����'h�ow]���$�=�.��k�i7�����e�-r�I�rv5���>���`|�B+dzV =(�b�
�B�g��$�K*:5:��V±���`�FjUْo�Wk�1+�689�D�>��c����f����8� �XC�"*�Xda��3�!�@/��U�;���j'5� U�ԗ	�FBq��o�C>M�����J�Z���0(F�0h7�*
��y���Lu��s�$}%�>�@�g{:��S�ҝ��^s�&�����*� ����E�Ah����.�tw�5:��]��kp�p	�P�y���oO�U���;��"(!�p�n~#���>��JcՔ-��YgNY�@�12���O��掭�c��m�Ɵ��?��C,�7��dގl��o�c�Y�3���,��lf�I�~ ���*9�{�Ee�Oш+�Cs}��$sGr@U[;��`~��qLvU�L%aH��aƀ�`�L�Mt�p�);> I�0F���$4��ܹ�k�t�
,~"��~8����M�ɩK A),-2o���zx���5=�b�^g��jeU�_{7�[/BJ��kqu��
ǯ��B�,���]c=������K�r��{�3���Eo竘����	_ M%@
��'[�ғz ��#\�|Cz!��� ǁ�޸����uYo[�����쳇�X���i�	�T�b�`��%a�Xj�gW��  �8:��d���҉��V @=�Z�4x��u��e��Y��ԥB����&v
ץ;�����N�U��2���^[��]}<D�}�|�i7*v�=Qw��<T�޸&��
]�4@P_���3;�h!z$�K���͈���{6r.#8�l��AqqB]h�1��^>0e�//E���rB�<�t�Q�N;?;�Ho�,��'��a���H(;t�Y�	�gS��n�<K	oV��S{1���N�X�O���%q�s׍L=�����U�{@��{nۘ���JgY�ُh���/��C�� r.�v�p��jdhEO6g�і������J�X�T�Kɗ��|��z�A�z�y~&16�{�f)��h����/��!úJ�L܉_�<�����wsJl\�r���i��Sq�wwgZ���b�|E$���������t���Vё�{G~��t��Jʿbd�k����4BtP��ͫ~벆��L^�� �du�R�1*�}�$f?`"J�.��3�.��Mx�|�}ƿHW!}��,�#�2�ت�� ���$t����L�4R��>f��,f-"�_ ~vۙi�_g#�O��}�������"�m� �Xq���q *�ߞzXD;�MO:��r)�pME�-�K�wv��@�4;�&�Xˇ����q�,fޟK���PeR�JGq�p�.k��q��i�*C�t�ѥ�����À������˸*�l��=�-c]T�_Eն�Lw��W��=�w1rFx�EaJS���� �,~<l^��/��d3)�C����O��(Y��9�`>d�Fז$@]\�#F#s�k��-��� k^/�Ğ	a�ru��DPB^�{��kt�[Դ���AQ��"֭��F:9K����;b����㬦|���" shN�	
�|К	>ɵ��;e:u/x� 1���fĔ�.����%�T��{�'�2D��
`�Ƶx�)���Q8,깘iQ�<'�ڮ���Y?��@7\�� )��xq���}{?n����Hz;��"Y����a@����O��1�
�"�Bbz�(!��N�b�7Κ#kVz\��N~�	�+���ӱ����yFT>����s�{��3-��q'��6�?1�v�b����.M���6�iXʤ�t���%�(�'*\@اC���1�.S;Zռ�XIEM��~�$ʵe�iҥ$�,^���j~(g�~ĥhR�3��$�窇
7_��j�c�lt��F7��OV��Z�������"i�"	�|7�XS��e9g�mv^3	�e%�:v��g�������f�U%�F��bY����A��n6�9��{�v#P�.O��E��);o	2��ݍ�;	Dp,Z��������c�Z0�\�Sx?�pK�j�Q-{�Z�  �!Vf�`���5�ģשS�'���}'=��0>��/j7���+�C�u�]�p��t�Z	-�'Y~��B\�x��F�T�|"gE[YE�Őy+S��ܪ�=��v��X:��FUݷ
����Ѹ�&��tXX�+��g�j��p�O� �5��*��N�����?;�W�UǶ�5g�`5O9�r�F�q@�������p&��3�����nq��;�;�/���V���_J6�<��a4�c�Q���_�g}���-��ހ��L��	O��.�׼k%iz�����������*f���I���]�*Ċ��5>X��_�G�0)�EE�,,.n�X�u(W�x��vO$aU���˪���H�;x�1�6
H*�����'��%"�;G��L���t���	�D"�[T�e�����w����̕;$��_K�*�s+�x�ל�)��r#�����Yh���ar^��#@�5�k���L�����X�ق����C��r0}��!Wl���r��Ճ�qM�'�h���$Թ"d{m��_�[Bt]7��H��H/B�-�6$��Q)e�}���ߛҷ `r�6�j��2�K�M��k��g�n��FU��	l�^�W�=��G������^��A�!ˎ�F0���&ɓ�J2�(�d9���59��u�p׿?�y����f�}��(rϠ7qϳ�|@�ว�G4��/Лقh~��4p�[�v��"~LZakTT��No��w��b6�lQ�{J�͛������p��UR��� �QY��p�,'%�{$�d.�����mE�} �U�\�7�.���1f`S_!���Hح�k�ë6�&'@����75��y~��%9u��e��I�D��]���i���Ȉ�  �"H�z"��M
��K���J�jt4R�N�*�yͩ�1���_g}N���4�z���!�>�v Ņ��g��u8jմ�:PK}��������l4T�$���I62��໠�yy�r��ם?�����.\�%�{�+>Z��獵!ڌG��4)����@�2����F��&��~����-�A�i�v
��n�v�l	6���,>.��=�:�i4,�G��}D�;��ۡv<�YZhq_@Z6U��k�0D ���4�y"8M�Ѵ.��%▞��\]!�,`��Ry|�<eg�sB��� Mr�c83� Dp55v?��Q>�$G��W �VW¹>��3���1{���S<��B��ʦv�|َ�7�d���P�[�!U����thE�|l�넲��`N�H>ҕpę���GG�.�v�7g��mw|�:��A��f�	ۤ؀ȞJ��;~�)���~�'�r<�kbil[�L�t-�<�&�8)�4z�x �|?T����Q|��Ut^q�[_	B���~�VG]�X��y�X��	����������!`E�}c�@
I>t��<�6�����h�A��;����.ِctS4��c"��W��a����Y�8s�z�2�Q@/JS����^�.�aZ�V	T1�'"�Uj��o�9��`$�~ޢ���#e�㮭���J�mPU@h��д�!}�L�~Pݷ؟}��=��:6���T"�� ����$���u��Y;\e'cފW�P�]��q׮�B>E�v�8h骩�O 0�]V>�T�C�2�g>U>G��Ȧ{�ky[ǯ(�O��w���^�p�:��-��Y���Ƭ��x�j�p�g[�.��J-�D���n��=�W�
�~fa�g��m�\����[	���p��֌�$����e4�T��É�~��QI�G��\K7
���dG���X:l��Qx�gK�ɐ'�V3g�)׷���~�C�c�Il�b����φ�v��`d�z�i�zR��s�+HXHf���|�q������Q���M��e�*t�F�d=�"!����F)�h3��yj��q#qՍ��JN��tɏ�R��(+��q�ܸV^w�	iK��:p�kpu4�ơj�~�J+�~�<��4|�M�Vn8Q���(%a�|X�_��w�ޒ�f� n�}������^�w�9Ɓl+�1��+�����m^�qN�+�Y�4~xd���M�_����-OZ�e���1�9f�'���r�i*3�T��]u��<�s�Tܽ�5*�}5��������ѝj�y�t�Op]��d��GCs�)٪�s�(�e�W��X/�O�5c�KR�^�w$hGMF�j��e�,��9�#���>E%��s���8�	��o��xLN$�'���YZ���52�t�GR
�7�J�r3���~oU������ϟ�%�7��1f�-K��������>q�?X��k���Q�Ą�'K��m.L�g���50�{p�IS�ʇ��d�5�ث�ͱ�;��`�+��)AXi���'�ׇ�������aX���؛3�K�@ ro���MX����fl�C��s-�+��؎<��!D!L��?�m��bS�	���W�AU#���ګ�gk>d��7{,�̐3=Y��{z��C>�����4{k�2���%@����lnB5 ԝ�_�a̍��v$VM��-�S**�Q��Q�g�mn�5�������� ���bb�nv`-���Y*���˄����~�n��TxHr'�-;f�-@x�Ǐt<���_V���k�	A��cl���C�x���.���NVUkj�5���wSx'������}�_�ˆ�~D*�����L�!8ձ���U����k��Ͻ��\�-׏�L��]�zjg����v���l%� �!4��c���Ҥ1�ol��o�K������&o��qGJ!P8�<���X���z�������q���.�oxKS�A4#h�[�7&��:=ݣ���z����O�Vds��a o�?L�� '2����B�ևrh��M��-���v�4����>ǌ1��L���Ng���M��1��F�J3l��c��e�Td�Je_H�7i�<aңA�=� 39E]Me�y�.@�i���r�N��C� �95:j�Ʀm�:D����Ԁ��?f�w�V 'sW�L�Vc�O1��>������G"�F��.�W��|R��)�gF7vr��YaH��M��Q
XlxV65EB    4663    1130{C�aZW?�����ީ�s��S��#���$8�e���������̕�)eсw�#��ɪoZ�z`�_����m�&��Bs�a3d��.�,��������f/5���ݙ�UmG���?�h�o�N�d�lw�i	�˂�]�f��hp"[E-(f0�X��yh���z�� t6��˅FA��Ei4���<M�v7�j��X�t��A	&X(��)�ۮ;�����Hh��r+������]B�A��\C��r`8��;<�$�� ���&�v��(S<���ջl�2�)��"��AJ$�T�*T:� *#�:����V�_7L)������8��q̞�pt��E��MX��|ڧr�H>�.
o�1;��?S8c9/�B��՝ë��t�9^�yǦù/��w'�o�
�c���6~+�nJ�RޕQ�D�I�	1�x9 y�?G��ǆ!~.j�y�&"���	��4Z��X�2���:0�zc�l]f��5�8�	��5B
M"��G(��6���ݬTb��ӳfm�"I�g�@�_��mjR�D˽N8_4�����R��>b}�@u>�
�<ɝ׺A�@k����B����n)�6��cP
����Qeay�2"My:����m@�I���\��LCӀ�� Y�hHN {g#�7+�=W���R��RR9!�d��lM��N��J��0�����})�
@����V6�������������gģ/��$C��j��k���>>�'��p� �?wv����~�avH���y�\��Tr]������{ �Ea��r���r�X(����^F=�/�#V���Nպ3*�K2�Hj�ͷQu��=�=�K�ܦ�b*�Q�(�Ab ������:Y�<�ԑ}�MP��L[*�)]�͍��	mk����B�g�`s�y��-x��Ub{��X_���[`	�;�a��R�R|�%��{eq�)hWY
D��8R����d�Ar��@i�_M�t�l�~rw�Z��F�'+� ��)O8�t���8�.��^5i����X�ZA�3��Ʈۙp[�qK53����L'D�WE6z�_�^��˚�f�5[����:���� �F(>�:7"�U������5�F���H~�6"{)*8��2�|�s>��7�r���oz�N��6D�#}3��R����F(X�f���@�C�;Z ����p��~M�p[��|�6&z���r�߳�@�ȗUv �߷.�[~��&������۫��U�1����P��f����� ���,��� ��u�nm9j��=#"�TҐ.9y�d���e]A��Fg�LQZ���񹪀�������|�o�TW�v��7�[U)T'�F�ُm�6]럠��(I��2E�F� �D���_�Y'�ƕ�e�����`��8��3�t:�������֤=)��hZ2��;���q2�g�����&F@B)��-���3#�qig_T
��NH�B�m=�v�����Z[�jN�/M�������oo�d!4uJ����]�W��p՝U��H�n��ʑ2bk%����)pM���|�L�l��6Nrd%7*�v��/��?�i�~�����N(�o����a�P93��M�]f����]����d�|4�Ƒ�TUS78�U�]΢�v��*�C6E|&���N�q�LJq�+�o���������n�E�{N��uQ��K��^ĎT�z�.T�10d�����
?]9�o4�a�����c������&b��1AV�'5?3�jzjc�u���u���$!3���7Ɯ��B��>
"G�)���U	y����v�U#�s��7��W׊�$�����_�Q)�k�?�u���RW�?m+���v2���'\��ã�C�`-�RN�l2Xv}_���ݣ��?���)�T0����O��b���|��Pt�b��y���ǵ�ڣ�� ��iq���a^*�lB�V����ك�����7%�/�7�u��S�G��_D�
�������D�������U��!�K���Jޤ�E|e��-b���jڰ]��-簉�+t��$#�؇'��8¯<������eghy?�����>;��h�����Ma�=�}��������ĳzrpF53g[�l/ �GX3��&o%Ѩ'�6���.qJ�h��,�& �NT�gW s�6h��MQ���Q].V=}�#�0��F��ŌZ>ܓ�!έ�!����*�䃣9�6Gi�7Zl��J�y����9�b^��?�@�hv�nbC����(�f\K7�udA��")_�د��Z��ޑ�t�w]��!`����:jx}1?>$������l�]�=��A��c����Y�U��;��?̡�2��q���d��_N7⎦V՗�[���I�ipaT4������F�TbO�R^�s��_=���KK��[Bc�����V�ƪ���Ҏ`vm2H��cCl+�yj�;0��"�q�
��P������҇I�ҍ^�f8"��L� {�"�3��G缡�9��2H�����s<��2�D���{���b&��� ��G��<��/��]ĉ=T/�)�Z�#�l��w�u���9<z�)ࡈ��.��~�3����:8�{^���!�gv�Ys^C#�lSR�N�v��~�!��6�,��jS	u�Ġ��ף��F��\ݵ6ۧR�6WĿ��3'��"��\�����J��'S�0�Z��2W�P���_��s�yʮ#	P�u����?��f���l����m��%�*�~�\p���������$���R�hJ��{�S\�w�ARy��I8cd���z|Vx<�X
Ϧ� ��ւHc���gzC�ך��;0���i�e��nB��tB���Y�����S�<��W���y-�-�0@5+�`�����%�x��q��#"��"9�\aD����L�dS�_�l/�����_�.;���}AXm ��~\�O���	z"�Pf��	��M�.����i�屟�d�e��D���|�*�?��!Y`=�MM������d��1R�i��|~»�r�109���w����̱�"Fp��'D�_\>����<,��Tñ%.K�q^a�*�8��j_g;B���;ms�+.��ɾ�/�1�琢)�l2�A�`�K�$�Ac`�C��b
�MZ�_���RA�(*���p��\�AK�\b;�0Q���w�;Y�VP��3סNGf*��`�_�
��z��N�'��� M���+�]"rC���ь�Èg9!H��$R
1�>�M8�˷�	ϣL�ʛ�A⡟�xA�-Ϫ��\���W`9��c��&V$��t���! �3e5�u; /l젶��Ѿ���~���򨫑lՍw��+Cw5��������v�����)��D���𔄨���w_��#{f��z�;�Aŵ���Nװ�TyJrJZ�)�yp�j��)_�8�"�rXDp�o���8:�.JkH��>`�Y�y^���O�U�6����� ��L˸$��R�+I%��H��\S���NL#�s;!�G��񊉂���
u"#��d鿮���0���p
���b�C�15~���x���ע��0s���a�Ev{E �;̖�߲�mݗ'����ߕH	�j�'���\Ѝ��%���7A�g0p
�J|+$�>'ꥋ~�JNM�d�%�_��w-�KQr��zVT�qi��Lܡ�	���%��9�N����E�ѷ�u�1�?���\=��P�e�L��r�U�"ީ|/0�\!�<��P��7��{�]Jx8�������!6(-�#�;�A}3��	�0�酙�/�4]��9c0�Twa��7B�C>����Гb|���N[�F���k��oQ��j���!�w�eJ@ص�c��������m���P�(g�C)��̬��(�vW�$u���Wzx�&�������~o������1����U�@'��R�Lz�:��,�B�S#�r�؎�3|�<��@�PNƓ?*y�����
���WJl���u�4�������*_`�<P�%�wE��KUE���Zȁ��q%��P�0'����-<���D�t
K�QJZ&<���>Z�l#@�0�ne~ApPOZ�u��:C�˨����俣7t�mo��5j������D-I��Zgv�ks��Ǡ��l��(4}fu� �����D��>{�4�oJ�O�'�I-iG�;�����&�6reM�W!M9yr�r��q�;z���W|�+g�g���{��g��Qp8t/c���ճUU�����T��v��(�z�`��D��������
 ����y{3d��7�����b��u���_���hb��_�wkAN	��P#R�r
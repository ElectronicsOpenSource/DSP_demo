XlxV65EB    21d9     b00���,St�/`�E1W�aN�J�e�X�ّ�;,&65)�e>��<"CH�ɸ�����\�/�W�ǂ�.���	K�]d[G˫��o���
���Ő�h��}�nS���ڋY��@��9-�U�3}g]��^G%=����L�Z=�(y���oo��-��mLj��M�^Z�B�B�_�����n��p,�<ߍ:�41�	y�H�
�=d(�
D���Hm0���VI�]������Y!�?,%���-���Ԧ����3��T���Wbd6�����t��E>H�R__Snj��
Vn��ƽ%����m�8��叭�B�i�A�ő�p��5 _�+
��z������c}�*�"�e�6Pt�X3���w����	>�c��)���ep؊6�/q�����i0wS{ѠP~��l�2���s��2����~�z��7^��N���,Gg�%����t�5H�a�n�8ޏ��i�f���.�.H�P�h8���l�<*�]�l�n��+��*�*��_1b��\��}�b��4}9yK�~i�
0^���F"2O�mt�w�M�7ŭ�_�}�K2R�=4i:'��Jۡ�v��N���ߞԏ".�iK㶾GR�D�1��S�Ϟ���$�]�9����ļ��C�C'�j��eVg��1d�h��p��:�ߏSt��y�Б
�����ʜ����9�|qz���I����bD�S<��p�`_�|h�k�9��e�lvU �xK�@q�v4L��m
t{~�#O9s�t#�ʇA@���c?߿�]��X洤o4�(�6yTI�z�d`Zi�����M��*�@������X�����$:�gNq�4%M�&�!u43�GW��H^����zPI��у�g�8��g�P8�8���{OA)I�Ytw�0rn��Rm��Ze5�Elv�4Pw��� .�P�|�����G�/z���lR�MΥ�`�`�6�VI�E+�DZ�75��2f%^aGH`(�<�0�7zz|U���kH7WP<�h��I;C��Vc2y^�#�]�w[;�t��m�3p֟L{��}�bö,q�a�����dP{���a F��`��\���ה�ȃ[O$��$ 1!O��]O<��V��7+h�%ؕ��H�& �)g��Q�p�DF�e�s�g��g#-�	�����4e�dMs����$Z5�=p����BH����'�4�Y�!/�(��"cK�@�؂��C����� .���oQ�s�J�e�Bi(�������Į��Z]r �b}_��>f�/@�5 ����?/p���_п�z������3
c��`l�����D�$���*���9���N��١|��[]�2�dr�L9���6��sï|z�q^�Ģy�&�|�_�	`ӟ�IKZzsg��δ��`�^@ƿO������NZ7/2~�C�h�͠Ux^h�C/!zf�[o�Oަ�Kv��p������/�;&rA�B�"�����U�� T=��g�0�C��W��0����c��� �[�����=+�S�{;
.9���D�iP/���O��c>ңF�`��L��{�Ćz�_'nG@.#�B�hG!z�"K!����HJBq8���y)FPR�ڎ���V��&�JIt{�L��a�[̨�Eژ[�D��jGO��'a������T�L0�u�j�q'��Ɵ���7���Z��X�P���(z�M���:S�T��T�C�B��w�$��@�DD�����D��r���#�=':,t�G��,�y�'=�xb�s�h�R}Zp���g9�~p^	�HAW�:��2%��{q�{ե?*����}o�?C��>�Yб�2��k,�:ip���4��74*������l.�U�0�9v��?�d�.}�X9}�i���(�LW �ǰ*�YV~�Oh�[Y0�{��/�k�dK�,�
_xBQ�+�~p�,�w��?v@�E#N��1�*��˹I��K�w�s��3E
K_m���&����\�D3U$T;�S��?~@zy}
��97��^���4K��D�n��pAd�&/EMRT��m�σ�*\Ѯ&���Q�N3UB[=Ȳ6C0󼁂��F�=�Zf�]��xyB�n6p�9w!�Q59�v{��
��K~�R"�0�����s�,����1�H|��p4��{�[�!�N��.��嵿�w�Ԍs�RE>�H"�|oz�ҩN�kB�[�����h���&�J�uAE�a{@�':�G��7[�����lQ�Z�y�=-!!$�y?��8�o�ґ��i��"��55]�O�9ِD>-��9�s����<�dP�!a�5�a	�S��@��g��A陪X"��h��D�@�o�F���]sr<~��lc�$~W�w�E~�g_��z�*���$�`��z�w���4`��xu�0��'���qC(E�����7����y��ΛG�-�7�9��Mvգ.����.GH:�"Ĩиōm�&~�QX�o�zX5�� ���SÐ��C.v�)��8�	=��+�ڐ��$�@h��ɫ�5��
�-�6�����7�&�u�@b�H��$�6��X�|H��?"P�p����1���V��)-~��Y�%jI ��R?��?�b;��a�qCVwm��Z���6�|�q_ ��0m�!��cIJQ=��s��a�ӫ�ƶ����"�>�tLx���>��v0��u�W.u�Y
ˢ��ہ�RmЇ'����n�l^�H=�lr���L����n��;�*���:h1m���&��gP�
�3T��޳[f���1u��v�
XlxV65EB    fa00    3110
Ӽ�f(����N����d3M��R�d͐if�=�܍�o�J���ɧ��>�k�Xgc���!Y΅�ܠ�'���G) U�����L�����5�Xd�2<T��l�d�B@�8�b��.¦���MR����Q��q�}4ҒC�H�E^���2`�4o��M���\g:l�Z�}Y��3���G]\��:@�Pq�cnoe���6��u���H�0
�ex�H��*��M��K*I=Hgc�ѥR���D���߷�2H��t��J ���~ZA�n&��LK �_JA
�!qꎊ	,QD1a����R���&m| d��|
�	����wQ:~�*:�?TGSZp��+��	�:�F�:���U�H��Ui���Rנ���)�@YF��m������?8O�R�j�,ïfJ�N	*����EE�SeXBux�EO<hld�h��w��.�i�{�i��,�R�;M��(�8�)�Sz�����ߌ��cO6:�a�?�v��%��Y��{W�(���S!)���!�"�O4	yO��K��e��M�p4~�����S;dO6~-t�eF~��h�v �녥��?���,�%s�J�$
V��H1\.Sa�$<{�>H����-�����z�ԡ3W1�;-�l���B3i̢�������� .�9[ʽ��k�� �(�9�Hԛ{�-��-eeb_p�l��%U�����4�L<��q���3*�p2�ح[8����
+��~�L��Ț��5\�:�X0F�����Xv����=Y���8<O�2�[�+�PЅt	�ѮW����fk����V�XSI&	�T���jS>xFC ���r���C�cp�8�y��V��-�%h�D�R��a�y��Z����)J�ŷ_7ٰ�|#��Q���|0�۬g=�P�N���Bg��VL�tL�%q.O]�
'�R.<>F@�R�H�m��e��G���#�N"y�p�sZ;,�˥0�-*n���A�����]D3<Z�3D6�X�bs���1a��yL8�%� ��n��ቐ+��a%/��4��qB����}�j`���t�R'M	�x�r����w��-<���8#0��_�������
�oj���	�d���VtXN����z��t�6¨�l��q���pqC�y �-ܱ��	�4n��b2�Մ[w�پ�"F�%�R���,6�f*�t��ā�-�X͛����P��3��2W��B%6���'�����!��#��ݭp/�O�޳�}7F���. �Вj˘���>e,�s&�聸�I�˓���Qk夶�&|7O�=���u��@>�CQ/��)-ܶ�%�;����:�ΧI��eX�.�1 =ŭ-� %��k����
��E�Ge�U؊ȝՖMJ��)�`������Ɔ��2�N�%U0hЇ��$�%:so���A�˹8��>��]=��V����\2omgFo�����&�e T�sF�ZB3@yM �o#_A01����{�E���Ϯ0���~���]�,U���0
Z��QA��e<�;*!j!�
��r���tQ$%#П�#+�H��!md���
�]����Ŕ�� �Ŏ:8�<7AP�h��T�P�A�>/i�0'��\���W{�D[tv���D�?}h����X�Sn��embw[ǣ��D�6�� �U��~�t�׀Y͢` �c��
�F�e�0��V]�"~f+W����K�� s��I����=�Q�EbT	o�.��0=^�"�1�p�a?�E�Z���>���tq����z�Sv1j��������s������P^�_N�ҽ����S�y������)�@ m���;HG��:�I�ˇXœ�'��� ���B���[w�t���4D�k�ճrr�ۗ�J��u5݅��q�h̾v2�{��z$k?��qh�E���k�&��x<�8r�E�Q�� 	B�1����E8�mJLpF���7|�[�(|S����C������T��_��no{�"n��"O*ܳ1	�DҜr�l�S6X�P�,��_{��H��W���)Q%���Y�<=U�Y�v�h�b}9��޺��e��oM�B�<���c*]�����������\�`���TQ{�)�M�OE��X�+$�gI��..�k��E�� X]8�����7;���D'O"k��s��B�&[Fb@!BO��q����58� p����G��i��n͋XʢD޼	�8���c�n�}"m��tMe��S	�8�K̭��þp;XX��#a�����_�f3�1���pr���w�h�����Ju���s�d��AS���8*�0�+����pn��y&s�qG��2�z��W^��Ts��8�<?v�u�����A�--.maz��{鱬����~�_ ��1R4A�1�+,\�u�G�g�N���hu��`���l��-q��	狋��<�/5�)Ȝ�ŭ���Q�m\j� 1.h/�'�Mr�ٗ���pە�ND�z�͛]4'9� �����?;\ωm���[��/ z�c�5J���茱�$qr��L'�i�!4��U>����o{�@$�Y��#�q�g��!��c<�`��������$T�S�GK���i��P��'Z"��a3�V�~H]�O�mu0�a�u	~�Fڊw��Gg徜�0{�c���#y�e��K���{�d`j-������w�o�`�������ݻ�=A�}�����G��H�8'z�M�2���g����n���j� ݤ���2Cxp9qcݠ�e�g)��le'������}C�J��Mz�O:�X�T_���V-�u�~ȷ�"��.ѷ�'/�kiX0��=>2^��഼��د��V�&���a1�z�=m�й���r7�xB�2��?����Ҝ�?���d�#���~8T��7�lM���pޮ��X`��I*�|�[Ϊ�lg�߁����մ��46xtX~j�'2{�Z79�=X�NO�;���%�WfI������K��s/@�|�^4�����:�-�c�#B�R�J����,<��=sH����@��S����vp������D���QS[�(6���ݘ��2J�AS����]��sD-������Ěw/�;�8+ݧa��:��1�l孡4	�{���'�\���V>.��1wōr�Aκx6~Sp>�ͪ�Q��,����'�.@�T+$|YV�!�G��.i�N=��,x���ѹX��2�e�a���6U�,��ԞS�r���:nḶ�Tc�oVo���m�/�̤Q�HZ������Ł5cbGPP9[��QDw��8Nd�+�?���_.���w�[��z���T,����z�@V���t���~j2�'
瞋j(�Lq���c|hk6�v0<����g�Έ'n?$�1v�}�����}%=�%G�4��Õ%�9�cE��o�<��[�=�ޙ ����w�b��OI�f�e',00Dx�L���z���hI_L�?@ �Z�V�j���(�/�P}
U���ep}�W#�4��F�-��Q��O�?Y�-��y����Pt-�PbB3�\[8+h"T�Z
�	热 �Ӕ?B�:��{N{7��ktD�Bf��UT��N ���	��S��x ��� ��SQ��f�S��P��η�fj>�V��d�X�pK�k�m\1���m��7bu���i�]⹷ �rC{�\�j8��oE��P�Fv̐ugG^v��`�����&�R�E�c@r���ub
d �P�I�ve��Y�2���|(�����8�E��":��$|Qe,|F[7=T}�G��S�em͎Ґ��\��cO�+.yE:7�LuQ�.��:4��a|$z+�+���ZJ���Ȍ�}��/̋מ�4=9sh$Du�h�-�B:�z��Z�qu���Y�]~"����-h����7�l�&�"�v���d&ML�?��o�c��{��k6����?,��J�86���*u��������SʟE�, �}��Fl��^��t ��JA]$�C�S��f���g-y�O -�_c�Y����i���F=/���O��B�����j����H�X�
}�2�	C�q��
IA��c����*&u1ձ�"������ C��rM�p�%r����Q�,A�D��P�u�AᜒűM�8�W
��t����XSY���~s|�P�)ʯ��A,sy��}핮�I~�}��b�*�p�3�T>�$�XJg�O��b)�3����� =�Y �*�R�ؑo�����q���z�d�7�P�4�@p"��`��K����Ļl�9D"ϑcM��s�N=�}�B��c���6�fQϓk��)������m�Ǚ�mo���p5>'��P7��n������4LN�qA���<�:��j��v��u��;~�S�u��
&��R����L2�^H�T�ilG���v8��Ze'n��̴��e��t�q�2dA�;�����x�?I��3���,�����Ps���x���Okg���-�2��x2�.0
 8k� ��K��w����{N��`!lϛ	7|+�;bU��_&�8�����_�=3&s���Y�3KK�\�=�)@TN:֤���f�l�%ڐ���U�1��S��{0=�p�y|.^/[#�Uc�>��uT�l���A��]����}�V�Ꮡ���j����û�H�u��(���{�%�P�k���
�%A��g��[�>�N8$�8�U#��b�t����gX�u1��F,�'G:`�'m�K��ac.s] ]�r���܁3��J��ZO������I�
�5����na9��&��3D��lKjQew�%�� �v�5�xD��a�����K�>�o�T`}^�� �6��*��Ⅿ���A�+�(�B���bxh<;/�W�8o�$���^#�Y�G&d��66piB|L��!X��s���
0�n�� T�F��۱L8C`�� ����_���4���A��b���1 ��&]�t%��ӷK�s
cjWx����,����N>�
aμ�/�9
Nf����,����P<�Y�k
�fnt\m�(�Pf��T�A�	���p���қD9�x>)W�A>!v*ˎ��L������$c�U�@>��Țc�{~�!SN��n�3�P�I�ȮB���S��N,��Ȉ��\�s?܉|@H��Hҋ�T>���nkR��6 qXu���Q&c�ҢM��a"%Ě���9��E^p��)�!���7��ޘ��Fz�S�<�l!j��~��@Np;�{�A�G�=Iׇ��������b�G̔!?U����%M.�K���Zё$�� �g�0�JZ�+�����yrJ��PL�YO<�I�r����`;�V��G������eH�3�٨�c�}���7���o@뒜vO1�K��ӅZz�iƬ�M�J�d���p��Φ�^���=l�+��'�M���;}��IԹ;$p�n��|�.'�l�`>6%�0D����q ���{�弒�X�|9n��ǎ8��
`*��У�+J�/�� �<Z�>�G����G5��<,XD,�e�$@T�K=C!��/A�d ��T����� ��@@�K��ʈ�2�u�\��F0o��#��o�\�����k� �y�m-?=���r?��kv��3�>�m_d�C<4�V(���&�'J�8!mژ�>�%�����V%߸��}y;�?C������lY%s�m	�0���j�y�N<p��r��cgy�O\�B	4�E B*�[��j�YX�q�+��9��Q�g�dj;|���&ĲK�I�W�U�q���V�2��[�ߝ�E����3�r:�����]Ix���K��X�y��w��")�^/+�E���^��q�\c�&�����dԃ�/��
΢�]6�XK�r�_��Y�.���&�L7��?��6̪��>X3�f��SJ
�����##Dg�o�Q�'��^%:��!���������A�ʤn���������m�p��a�9%�$RY=����1�ŃFtU�+x��T�5Ú����� ����-�AvZZD�+3�����fk����Ť ��6j�%� yt�'0��Q�`�b[f�{���x�f���>үLňJ�kq�(�����X������O�
u����Yg;�[����ql�M�[v�9tr�s�#h���^A4	�;�\��
f�Q*jjb���w�� �M��Ϥ~�"�7(��<�+`nt	58�yWQ����Ul\�͠�L���`�pn[������.M���������_�iaЕ��p�Ͻ���\n�/��vݷ��4�X��=��P����f_�,OQ�UK�_�@�y�'���䘼P��(8�$�	��U�`Q\��Qza�jE����#Q��qs�n�Dk�X�+�o,
q���i�:��\
wh'�b)t�x��mA'wW�]T�Ca= ��{���i��L��{�o�Lm�/4�ϦK�e�)å�ȋj����������:�6�#A�90> ��g`ً��j)�0���F9�b'Ag��#�W��E��ک�[|mSź��[�QC�f�Z�6�Q�XW��ۈ2͆!�D�9G�T�S�nhvR/���(ݚ�e/׼�q�Y��^;f�K�/ZLŌ��[�x��v\d���;"^��:M4�w����c2�$m��[�7���u&����8(ߣU��#l��E�5�OF�xA���mpm�pv�f��u/�6�k��O��B���~'U��bh��V��6d�&�W�1��
�D��!��U�Ox�� P{��@�d����8��ȡ?���&H��{�wB4�%߬���WM����Z��}���O���%�c\̌��N��Т��Z��m�I�I��� !W1R;LW�i~q��e����աY0��=�R�Pߌt���ҭ�:L��F��*؞^��L4_�O�����߅3�ݣ`�܍䥶���:=��6�{�y�g� ������������ܢ���3�U�s�\1���5����y��1�؇���H�a}A�$��0���=�"�Ds��G�̺#��������
=����ٷ:S�,!:l��Km����zq��=@2�uˠ��<*o��L��7<�c7Hޤ��/�C�!�)a�S�~V��RpC�m�8aO-�5�Zd%L"͡��p�=���)Rf��,�o�Ə��,µ
�-�J;��N�5�����6�I��pP!-%�BjI"�z��F�m�,9-��t�7Vʩƈ :�2ym���U�Z�P�`:�jcV�狾�]�x�Jx�n������D0J�*��Ǌ�a^��R�پ	����-I
k� 4T"��~�/!�׫��]C��; XP:���'vA�4��Н p�����o�">����Q,'r�ȟ�Zʥ�I�N�V~��!t�H�k�ZP�(Wcyi���ذ8����KJ���`@�Ӎ�_��R��HӨ����L_������e^8	��Ǥ��d����*��ʺ���^T���~��BH,r�
����8�즮B�7����T'������Z�w'	M�P����K�9��І]��
���5��A�Ψ��o_�D���@.����v�x#�F���,!Ɔ�qN�������<].k(�Q��^'�P�y�#�R}��m7G��y�"�8o�l����G0���ҳ]$���b� �p�0B���Wi�ޅS�{+��q�� �+ӞP��T;/���w|��*�&C&�o��K(J��L1n3ʚ���Ԅ|���-�_ċ�4��
ꖦ�r��?\'�n����M�OlA� ��2���d�E�\˥��mD-��m�1�GD��$u�_�B�z����G�-o(��{&	$k�)�w �QMu¢?�A�O"zr��
��.�=�Yʌ�|7~�(-�
�{���&X��ٕLm��'���K7��dvlvR�#_�o�W�W]��=*����C���3��mǿLjr�>�b�r�`'�?�9��>j}���ep>m��p�Dd���0Pm~[�����@5�<�
Y^5t�hRZ�%���Ư.�yE} � �d^v�Վ����V�u�;��+M��x��aH��kh'�y���O)h�OB-��M1�Lǫ��w�vkf�p3���"��Л�r�oa'A�m�kfX�Qa��	K�ӟ#S�Bn�k�4�G{I|��9뎐��敎mY] 6��{�j�R7�v�&_L����W�6�,MO�t%}���a\��R��I�V����4�2��/��(wl�mR�՜�#��b>�~Ӎ,�..3�&��sT��Lg�G�5n}�n]̤]�m��gU'V�l@s:���J��; �|vǧ�pұ�+ F�S����-���[�Q����OBZ����4�ɖ����1 {(�!1 9�R(��-�� ��	�W�~\�'�2�w�#<�ծ�Y������9���n=���?O�N������ҍ�T�k���*O�U�Y��5r������3^}�cUR@�е���2�E@VH�!Vp����#CbL�����B���8�%*��=��$�!����:qv#I%
�~����(�x� ���%r7L����Բ�RF�곈gc�7S��_�56NxV�M�)_���1릸
n�\֡��ѣfRo��6'
=U�T�w��c_��
�W��1�꣹�S�O���-�w �\]�N�s�6N�� �T�O��M]�@�$wl1�d�l��p�1�2��6ɹ
b2��_3�D�	���s�8b������0����bo�3]�wN:��n�/������m\��yY�VS��~$������jꋾ���piw*���g��%[p��l����s��#Uz�r���ԓ�s��
{D%�~
A���`��[��o,O�_��yl���5��e,�A�h �m�1�ocg�(��1�{�g|�^�^8c��q�R��f�K'��v�A�6�rУV5
a�� D��ɼE<��vn'�֥\����`�`��$�ޗ���q�����~6�x�Ʋ�t(��u��-Q�1���K?g�0=��꩷
���U$�m����
�H��/��J�7׿�x���z4��c��'>b,�O�.1�Pʼ�9������],s8NJde�:��v1��`>��IM���YB�ag�ջ%�`��ؒ��b��[��([W�J*Y��������x�}�8����W��Rt���fy���џ�u��������_}Ysb�Ӽ[J	�[�}&L��@�p�Y���7p�~5��"��k!���Q��6���r��ˀ�D���f��)"�n�HȟL�22�i���"3���2��^�k���.��7�\~W6�^"<J��	k��Xx~-���,��ԹQ�����*2>���Bӡ�!v���&����^J,���Ϗs����oN0��idې˼���&��"uH�5�t�4���6|�蚘[!��/RP+2)!�`�����V&WNR2(�Za�L�o�_���Z1����J\VKJ[9�����Rβb)�&_�9������0J�0��i2G3$��,i�Ǐ>�3%��=P� x����醧XM��v��@��5_*�a����c�M�AUt��\x�P;RϤ<9SQ�4�ö;a��D�N#kǢ#;��['�`��$�8:�o~��f�§p���j��`߉]�<����L���s͕�l����@Þ�����L.i�K~ٚ��h4�U!�ԑ��x�1�z/�W!���#c�g�㙖��ÿ�y��+�~��G���@ggJ�;��s����C����ϟ�b��� �Ш����D+���ǳ��5-w��O��v2�r���ݏv��Y�P�M��7u&��lFu0��h�f��I��]\%���y�R�kϪa_A<������j���c����
�S��`�5G����H��J�,{%;�y� Y<��Pn�tdcMZ���H@�RI� ��Ζ��*6�GeS�.Q�����s��`$�^��f��H�_���. ��c��6ţ0֘n��K��`��w��h�g4�3v��%��߻��
7u��P�w⅊H��.sܩa���g�l��dbPY5�5	�6b����"^"J�Dn�M&�������n1�i�����x�5�N~L�h���	�hm��8�R�`GU9���Qu�t:�e�Q9$��@�Y��P|uQB�p�'�г�U���Q�Y[Z��O?2IK�E�4��ɛ��Ldm�jΘ����a��$}͋�Y^=����$M��5�o���Y͚�z�(2�Te�w���0Õ��7{+5����K/,L��6��N�q���RT1��m�,7�T���{�zn�t�u���G�UǊEb7iS!�� ΃�ʪX���̜*YU�9(�G�-����X��,�=�4��JL0�����_%��t�������~�̛�h�-�'�#�K�עh_�6�tm�e7k�����H1��o[~��U���%�Zoe�,l�;�ֹ����fw�39��t� b�0Ym4iZT?�Ji*�#�S�eښC.{��qLXh���k�"Y�p�Jɱ��po<[�����]���;O��6@��@r�bb+cU?X���:�����qq�c�g��ҕ��ZV�]���)H�33C>��*�t�^�������\�6�ÐM{�\X����*� �7�p
��ޱ�3�5�^�b]�qJ�&	:Z�-�3&>˙�L�݆3�%�'��.���������}��;�<�kc������24�� P�OJ~P]�	N ��#���wS���§qÞ�a�w��:�>����g�+&���{/㐋�ɛ[�A�x�3_�\�9�E��P�`?���ly�v��5Ｂ�('�nԌ����K_�O�I�HyoB��	���_^+�JM�.l��E����um��9#����~!��"^�y �yU�Vѻ�N�,wC~W��^�:�@H��]��3��Υ��r�2WR����ٞSˊe/s�W8~���R#��PȎ%F�ϓ.���~�����8�3H���X�o��jUٟE�u�0O!�U�ZM�/��},���q�3�M6gׁP'�=C�LI��"��'�3��)�83ea�?�W����?;����-
.�	T�0.2[)B��Z�����к��d
�z����اA[?�d�-�\�N�,1���5qYJ9"92[���aPk�t�S�L �+��Ę�V����=�-��Ͽ�Q��}&��
�� [�u�U1E;���9UYM�!=q�`N[�t��]i�@��s�x\^���V[H�Y��5�bx�<C���^e���r�j��K7Y�v�`����:�� ���t��͵� ����*�R���MG'֏���z��oF	���!!S_
	N����^|�w������W���=
<�l�d
�3}׼�{����CS]8������f��v�����BP��V��}^=]�K�(.P���n�+w�n��Z�G�t�}�G�$-iK;5/�qKgҕd0eA�6 ��'�`]�q5��
햠kLH���<62�O�5O��o'�a�6�KnYܰ�1�� @{�� �E�h>u�E�cx��M�V�0��\��r�%7�Mi���s�O#I�_��L8�V�V$�jE�uQ|XY�~�2Z����R��`ge�|��F	:���z���#����e��Df��#���z]
��b��:���/ �çʁ�W�I�g�L�V%<Ws���Zo�%&L�| I�R�h�}=�r�y�</�X0E�NVa��{C�bTb5t��6	�Q �Ns�x�ń�j�H�
����54��S���a¯��*}����A7O�hbB�!0��2��R���k����. �7S� �iՋ�%�������@'�+���3l�M�N��5�n���ݍ�h|��1k��T/���>��~�ds�+�/�g���,�7E��1��Ʃ/���n�Q�U��I�.N�*=�w��m:N��3�-4�R�������e��4��
PD&Q\<�T��?*6�\��H:0lt|�����w�'M��;����w�-�V�ۯK��6�t�&�^�J���	.,�<s�wP(�d��1�^�ۋ����K�� ��op�q�����!E]�����1��Ǉ��c�]ⰧM�4���n����X/	�p,E�Q ��F�]O��:�u��'��}�V����YI!�y����e�2��)���|cf�I���
��Dy�щp��g�Rˍ�x��\������-��Q��P�5y�q|9����i>0��B5���;
]ݦ(@
��E�5PUR+���<�ɀ�g���ClXlxV65EB    634e    1230ұ���x�o,^�(��*Vi�Hs���IT�����L@�^�����r6��x7S��	d��+e���K��.���G��A' Z�"d�z��K��oK]�N,�v����#�ۙ�뉔Omߡ�e�-�����9�0f��e0Z���c ���$�1�[�C�`x�`灂��5A[�-��c�N�������v�XZkˠ�r��Y�i��u~��H�v�Ū��;�����p�}^�P21�(Hþj��ԋ���L�"%��>U	y�Z�xV�����M	�\ɋRN4������� �w�qK�(���]�?5N���#&�bms���Ci3�s|T�D����;�K����į �rW��\�<ܲ�iF��D����.3�6�{2= (xWKNjD�
6���	<����ԥ�q����V��J��8A>�[��/09{��n�ehV�vcy��eE�
mUJ�+���K�� ���H�r����U?�;R
�{ay��U�XubH
f:�Y@��߮p�0�?E�d*!T|��W�ɸu��Sx�~W����D�0�ؼ�Pim��S#�I;G�d�Q�����G؞�T�i�nV9~:�f�
B>�KmW�IS�#�Û��^�%�]��}�I8gcN�MB�(�A���W5�@4x�5���+1!M��Lǁ^�B����h���1���E\��<�G�l���/�ʇ>�ڱBeu����Rf�U�Z��#�/l���]�����c2����p���wi�w��=���fw}�"��E���HLG���W#�R���/�>��#�edAf)-v�6m��[��~Z���?��9�o�ٜk�#|���2�Bj\H�x�T���c��U6�1tK��:����"Ʋ��ci�e*�a���tZ�bb-��*��Ec/>�lGp�冠���;�\��bX�Zv&�H��C�n�"4C,`�u?�ԝ�aiޯ�ho�D 4j&�dXVWX�c�=D� ��Lһ��hs��Pj�ބ�w��p�X���L()�.��3T�֚���`�����1UOl��������ϟC���"�uP����<-�R}=�Y^��(�lk�z���������Z]�=�uw:}O���k}�`���4�q��f�`ke�d��ztb`cǧ\7��zn�l���O������z���z��?�T	���p"
sÄ­:�wd�bg81����
&�w]x�L�����Kz�%~D����"�6���Y�������4
h5l��v�n8���t�<���1a�=@'��3�f+����VV��ͻ~�<D)�z"b�N:�$�Ă�W/,�[�}�f��t�^&:�E}aa~Y�枧p%PVV:��5c�\=k��
!L|��Fd5��v���k8 �dr��+V9�QZ7L���s�������;�����h<m�e�:#�/�]՚y��H3�h��L=I"[��:/���xoC#�\���\ɿx����q�T9 ����f{�I�r7A�	�� �k˩����|�S�$���m�����+�ߘ�q)��rc��l��:�#��F1�%�:ճ­Nˁ���d���nU$�/���b��̄ҟ=<�[�kʕ�
��f�_�!{r�l=����rW�n]�l�f�rr�2{���c�2�]{���5��Now��������£²+�d��� M�4�2d�Иc���}ǃ���[��-�,O�z��A�`�TX�;����h��G�]���o+�\ �2��Ŭ��Ȓ�r��0%M{�$릚��u������2k�R��8Y�A�?��O�p�/�%r��r#��S�1J�o�+�S�`/�H�#�vȣ_�z��T��F�i���~uJ��2�7.)p�S��缢K��m�h�c����.H�����~��1�Ǻ�N�����_ ���
#=7���;�ف�sV��O��h�	���K���ًͽ�	�+�n��Á���a��Q+I[/��aH�&�����99/�߱7[?�9~�����������Y@_x�&@1�Y��EY���A�aܷ�?,"A\�!�|V:���	󻫤���wz��0��A�x����8x��Y8G�0y!"�؃x��I���VGd	�;5�
�E��a��/j�����*/G��>�^o��? �e�:�����2��v*�@TR�Ͱ2�T}5�r�z�p#*2�,��R5N)�M�����E��F�򰜃�i��4�4Q�����Y)iql`�����wv�h������s�ɸ�c�-H�Mw㸣Ջ]���&��g͍��4T�>X"��h�toV&]j���\o��J�=�!�5���R��@� �E��BR�I��x����o�,>>C�I[����!�6N�6����{��F[��Н�s��N�Dt�
�T��3�}}��;��x�g@��h�Ͽr��R&Z�t��Y�� \K+���!�l:��ɘk���xr!U�U���9�!pP
2}�h��%��ZF˖�M]	@H%B��]R�9b�z��� �V,�W�-�2�A1���Qs~	�uM"�p�9����xL��-Yrn�/e���4psq!Z���܂�>h
�K��S���9Udm�|0s�±}u���@C7�f����0h�4��Q�j�IbH�����K���U�ü�:T��(�aQ}�f؇ZU�Y-�������I<������I�i.Ls�`8�'�E�^K\��H=T�
�N������j���{�pkO
��:��}��p���D���m�w�Q�7�LO�|��I��X�,y�v�S�Ն�A��og�@z����}�6�Z��
&,��N߇y@�Ћ\�G3a��"I��",XǟTX/�~ȅ��s��y M�?��d�J�5�Mu���Z��J�J�aii�u��O�86}9�[�gu¢ao�혐Ja��j�����R����O�C:�Pt�����R̲�@#�4����vd��W�'�m��xu����ն���Z���f��D��:~{�zyt�1��[:e#��n�S�bv�pn^cg�s^�ʄ�H��^�����IA��z�\�D���+��p�-�݄a�-�A�r���@U��Lt�y��A\7vJ76���9�DL�+�B�:qC�H3�Fj!@��K^>��°p��\D�SH6��-|D(:n | �3w��j�![�Z��z�����b�b��#I�+�;)!���Zz���}���XY���Xz7�ă�3��ysa>�:H �`u)�_��O���`�sl����~�����+�A�wTm�du}�tx�M�6�]��؅'	��&�L��SM~�|���#}UM����L���'�@��1�"X�V�"��lhO�r`��e�^r~�!�j�q�t:��s!*��9^`��f���16��H�ӭG��Z';FҖ�Ïh����H���H�=��� ����N�|��	����x��Pn�ּ��7��z�R,h�5�E�6�]��H��|scCX��qS�K@JA6�\����
f>�-G9�w.�A�>��A�ˋ�iಐl���KI��}0w6w��W)�s�,Y�w`?~�����Z�~��OVS��<��*����<�5N��J0�!��e<z�se�(�T�!!��]�fXU;���&�2��.fhᦕ�Wc�l��h%� A�Ugt2�n��"C��ۤ�7n�)���f�-AB' �����p2�������������>o�cc�_GӝY=��b��Z�o�~�����*����A���c)���^�Ն��/=����i�ZBlb���1�-� L���t��m�Q����8�p	���=s�r�P�q_I2z�*�a�`���qz6��kK�{��;�Ui�qzG����P�ΐ/R�!3�	�O˟����8�,��֨H{ ��n�Rq4N�m�Ci&a澈t��!X
�%�'��*gn<Oq�d��/���x@h|�s��x1�%⮨qe$��#�wt�,=Zy4�A����뺎�S�j�����`��`P\E�������bL~�bI�1e��ͳ �k�P��c�@�o8��;����	�g" W&�q���M��������s���9ħ,x��Gz�Ft�U(����"aMTz��2��A�E�vx��g�fP�̖�5��O�VO�pNߥ�$��m�Υ4��+ƗM�h��3vq�V������g���vY����G�̤�Z�R�6�j'��}ձ�i��Ms�(5b�-+������M��DZq;�a��ρ�l�yOĳ�/�������_�;IB�r�T�}�olJ^���Lr;��@r�R4�G1�{3�_<{������9�g��xZ��-��7�6���(u#����� {���`�t�
L.l%c��y��s�D2p^��I+�~y�~��;V�_4��݅��K��R��G�9 �N`"ܢ��:�}F�-G�k��\���ĳ�xh!<���Б�!���ֆ9�k#[y;2˩ �6�?�2H��9������������T�H��"��J��]�6��Ͳ�3�q�HL�<Q#O��7�TJY���~E�[�
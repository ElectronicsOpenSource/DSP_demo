XlxV65EB    fa00    2a20v��f�(ml2{�lއR��5h�%R��T�0�S��>s)�׎ǎ�	�-f[�Qe����$�ip�f:��(f���C����X���م)vqu�æ��0R���ۚp���
+��ZzS�a��$r�c���� �E��r�����1�n
�&u��-������=�����QŶ�H��o�G�E*���g-�<�^�q�Y�����Y&sK�θ���V���{�XrȨ���v��B�,�O��2
�1�m�=�cE�Tɯ�	+��	��Ѵc�X�	q,�M�h˽���!��mK�L=6�eҵX�	����q�U��>�a����۰y�o�|��2M����:�O\����-�ۖ�t��v��~���Gb �l�-���lӯ�9�bB���p��������	����v��kr��*]"Gc�-��MȳY����q��f?���qK�1���7�tޓ�GQ}5��3����l� �kG`^)Q}{�ďܪ��wZd��'�O��mwZ|�9�g��Q"�AO ���SM>f�OJ4��1/�+�s�@zj��_��M�U�[��b&�� ���\�@����I}�cE�-n��z��9SB��8��6�vL"Sn�:)�M�u���)�_�>C�灉��sl��������5>�G���Km�����C��������B�^�Vч�}�!B-A٤�p�gvs?�A��� ܂�(r�0���4̭4�9ʛ��L^�*�\:��'M|�u��������;�0;��7U����h?j�9Z��A7`��a���=G�h&�����
��j�ġq�G��y�mַ���
�!�s��<k�n��l�p\/���ޛBW��̛K��Y�Ť��D��q�#��5L.~�I�T6D�{sK\n�L��Ŋ [�!V^B�oC�����n�񅒸(Vr��﩮�ٙgu�ݩ%�e���8%�f���E�|�;�*�7Z3*��D/6���g�g�tm��l�l��<�~T=_���x[�,�0P����'-K���b�q�5�$lh��4��e�VK�� ���9(ybt���A7v��zJ���� S�v�y��R�g�O��#-p;3:F8�rt=*CN>n@MY;�l�b㸘�5��σ\�(¤"��_�Z�6 ��b=���J+�[T|�z���0�t��1��GZ��4� �1�l[�Z2�Dz;ɉ�4Z��Fx�f����;���w���S�z��B��a؄Np�7��}N�e�ȓn,��t���/AH�%;��a�%#M��S��lX�[)-��m�p|4��%ժ�=g��;P
�B��e���#Ǌ3��8�u��cӞ�i����(�m.���Eq�VMEuuv�_?󅐩
T9�����T���j�1).��ܔ8�,x)����͓����!7����vd���Qu�Ά��U�_V����Y���P; &�/��ql��/Yg�4ʟ�Lx�u3$�)�;��|B�l0s�^�mANɗ?�vձ������1���.�_i��֕���-�R5�=-mC��IX��"��߈��Xx�w�&O��q'c%���[��L�ur&��������FZ��P��*�i�}�ƅ�@.��{�s1�U�h���L�� ���5��p��l7GmүF)ȧ�嶻�:IX?-���t6L������l��SF~R=�����ǿ�D�m��秗��N"���=,���������1�$X���FV\�l���16"H�ݩ72�� If.�S��lua�Bq����_�����Y�o_q��Ѧ���>jL��$Ri�Kt�����(�
�������~�%��5���AB
QQR
����Ë���4��c���3.���tT#䬀�<}���R��B��yèo��x���X���øC[�"�3�Gd�l��w�8�g^��C8ze��_�ÏӖ��G�ttlr�6TTA�@k�|+5��� ����N|a
A���%�@í��K�L+p�.�	�sS��y'`j��-�ͷ'��9�]W_{�d`A|��Y�x�e�xev�?�}ƺ�G�N�U	�<Q�.��l�������qe-��
�$��=k��2d�;vTF�O{Nq)��"!�<���w�GI�w;��2����s�����e��4�'S�$�x+�/7Ǒ�yO�M;i: ��wD�Vo�Cn�hmcE�t�L��&h���Ò�8����6گ�#����k��q���4BK3�J����=����-����y*�pa�1Z®�t�<ޙY��a۟�AX����qm�P��SY2���?�,��Z���e��0�7���[ZА��g���IR �����(���N	��t���=/Μb������sC�����G�� <C�w<Õ�yx��=۟�܊�4>�^\բ:��^U⾭<cd
U����O�`V\���B����G`W�	�|��{�}8T)Q
m�s�n2��7I���p%�8�"R7�x4�O,:���11|�>忦�|���.���#C ��)e�W���n����n�B!�]�g�O9�_O3s�Fޫ��e���%4��:��Y���."~�����r����:��w[��Rt�9����vP_>��f�K���z�ݽxLh�7��������PP;�q��>H%���m�V��[��%!�L�x���<�7n��3����U3�L:���ťEJH��U�*8����0��fy,%�.t-���r�<����g��l�⊫����ܾ�H�l���a'i��n��&$M�wF֊�m��֢ޟ`�ui��%hԃh3Ou��L��{p��A��]��Ӊ7d?�A����8R�ͯ �����t3�f-�}��Ve��^i�ȁ�e:BE�
�6���Vo�M�%����
sl�nW��v���u^&��%f@SR�I�sa��vŤ�l������t�k�y ����y�w������N���b׫�&k+&OG�@��ulG�M��i�u��ڴ��R6�V�7V���$p�[��#J݂�!�ȿw�������Ĩ��Bt�6�k���T���W�g_kPД��.�~���%�����[h�xZ*)'�'E�#(��9+�\�%���L� �xv����ʘ>��\]���Ҩ��L[j���I�M9Kq�my�S���2�{xA>�C��R�I���_[ ����^��])��" ���2} !����v���=�sy��X��������:���S�-���~��M��l[�L^W��fk��|�	8���l��nY�
'w�?�T�Ծ�Dn-�=�7O+ܧX/��vvd�����D~��)ptvZ��@���L�!>�I52F|���ڣNN������VIu�g6��6���0~�X�Ĺ�{��&^�7��Zď2N���;;��q�����ܪj�S�O|�3@�M~�k]�oҵ����T�|�����a�g�BBOD�!��$���.�@�)[~�Y�n ��[�6�~�Zrü�5�
����M�$W�K�d��. �Ry̗�v�����:��;�G�e�׆���PJ�a�����`{3A�����ot�|E+��ὔ3�.e�������w�W#�q��)�ܬ,�mωv�/�. ��{��1��|	����s9��jD����Y��s����+�{�4_Е�����b�熞Vb�1���c��خ�K�KQ#֦Õ���60�Rɝ܌*4��x͗��Q��`���=��FT@�v�u�|,�[ʥ��M=O����Y��N�����_��I�%Mr�"qL���k?�U'�#,j�:[YoF"$D�`m&������s�)p�*/aܷ|u-�v1V��KK �/	�bX�/�V����S9��ƌ��.�Q2|g�<�������\ڶ̗����1���t�7�]㨯�m��#>�GQ/���!��2�Q�������%h���_����%���ԕ���:��ޒ.�ϥ�,�t�vD)bkr�UQ,�Qpp���U��qQr61�V�('}Sz��{W�]<Y1 D���w!��G ߿YV�/X�������g%��V�K�c���z�vFBǩ���D�j�~��P�5Fp솛i�f�����5k�1�v"A� hV�K6���]�1�g]4��@�3Z�[l�d{v��!�A�T��m�� ��^���f��n(R�E��&?T  �_��`)�`�sc�Z��#O��<�ӛ�j��"��;�HE����%�ϭ�5s%�?�����k��1�;-�i����'���lqԓ��r�f;�����Ҝ��^�������WRh�anj�rW�� ���F���G�J׻�����3���$���%+����Q�r{X
.��5�}O��7l��<l1,��5�?7z�S��Ux���6��P�?�T�Hl-��$b�G�3Q�q�vt4E=!Z�*�k�n$��!1��+��H�Y�K6�^��%(K�HB��􌓱�t)�U`�7�2�#��49�)��gS��s��y8�%/��J�.'�@��]>����@L��>�We�yfQ����u�&�Y<:��t-ؽ�(琴b�cD7p;����B��%}��t��qa{�T+c֓���K�\h3S��HtIf��������ry@e�ج��K,�GC6�R��c}�]7w(�{\N#��l�?e?^������3^V�	_�9"��t��=�;�4���ks��h?�ˡ�=�3���|5�*Gx��5v�[��x��[�^B�� ��f΋P	b�s�
��I���q���jp&��1�*�ݥsG���d��¸����*`:cQ�g�� ���	:f�D��K(�
�V��h/�i��j��b7�p ���>kl�';mH>G�T(���{d.1�a�����saߛ3��U<	��0��C���b
~m��OT��^�&�Ɨ�i��)'�YD=0�E揬廨L��U�=oTH�p�{]!���w�K~7��P���M���|,X�������{��pVA_���[�9�Y�n�VrB��$L~o8���Q�J6��(�&�f0����v��څ79ؙ;	h�a��ّf�Z����	����1�	`��ȣl��TߌC/���7+���v���P��'��p���,�ra�m$�~~�Tv������p�	i�"��eD���t�=��΅�)�kmN���9k�h	m����A���[y�2fM�M�0�t,����B�1?B\���9S�7�ZY��߈���ٿW)�^�����:%� s 5��� b��U�V[L�=��A��s��e�qP�J��u��xjWR�H%AC�}&Ă�"�������W�Q/4c�cp�R�\�~;�&���hܩ�t��:l��j@'��mr����������g#��!{��Zc����y��L�\-�IW([�m�Ky;��fXA�/pOhݝ�c��Lx��o~j�2-4h��O���3�ͥ���I<�����,Y�O��4�ha���8���f_iYS��v�	:1���u�
�I�y��C%�������R�l4=g����kh?����e�hU���	��.�����������\�
�1#��#5;�s�����kw�$&`���7{�<r�ws*��s^l�>�%��uxj�Ho���}W�V��*K��W	�T����E�U���w�~m\���1�ozL����U6Y�?�)�ja�q�A�f�QZa�X0!�����Ǫ(ܶ9��X���O�E�9�zsѰ�ç~⣭L�Mj�(��]B7�R�OI��+����8��^�������r�J�X ��[�ʞ��b��.w���n�~�����gh�(NN����7UJ}'j�HY(̫e�[-���
�QR���f��*_�k�j}?pG�F��9��I�.�Au��mZ��sS#vl�r�}v��n�Ϭfc�߽4x,�糺Q�ݯu�6ԧ6�$�N���̺#�})7T H�9D"��.)-oJYqu�'��z���³�G��P&�t��+/��؏O�����9����k�l��+h��պ�D8}*`��D��t�u�Dr D�H�4/:���E�
C�;��k�0�_�u�Q���׿Y��@��4?rձ��-���R+y�љ�zMSqR	|Ks��5�n�t��7������t¸{[g��
����;����7J#d�I�6��- �aM�ش�վ�t�z�6'	ۑI4�-7Seh���^���*���`H�<�.Z�v�>]k�����"U[?Dd7�UelG��(��C,x��G}����YůA+�S4��'����-eH�����Z�k6-7)0��K�S����\ ��1�'j�	ؿ	�����6:�l�+�����C��t5N(>�`]��2>!��˞�4j���Pz�8f�m*�5�Od�52�����K����	Z΅��\;d��c,pX��[]������f�F����HWJëȲ[�(W��h]9{Igr�女�?�ic��h��O]&δ���E�%���֭ZU\X
ڰ��K+�����������㒱d#�tv
 Ԋ��� d��q���oL�;���2��	I��H0�����f	܊�D��t��k���h�##)�p�_ޛ�9Š�M�]�k.��H�׈/Xniq���q���[�U��g�:�65��6�.�b����U~�>�L.�)��@��$���y$&�C4i���Q��qę�g�?�z��c�b�٤��sͮ��l�����Ε[{-^�mT��7���MBf�l82���|����<CHMO����Gra7&)��"X,P�>�v�O{�>�D�!��/����(�V9��Rn�foőGϦJ쇇6�.�Ո�����\ZG���<.��w�)�rS�igqU�]Y�f)���A�-��,�TJ�3�Ia|xyH�x]N)��m' y5ɉ"~X�K�W���}7(��5��UN^`�bݓJ����>�~n�٤�Y������y'f����6^a�e��Li6����(4H)�-2�U��8�M�D��>���.4�o	3��=ř��x���"�OY�-�E <k�d���.yZP������Cl����&��G I��4�#�^u|�����=�#9ȯ��p�ص��j87i��9���ߺ!1�n�ݵp�k�5D[ W1f�)��{L������-b���/�:�X�Bp,�ch�jIs�a)ͣޜ��h�\�a�G�/�Ʒ�>k3��=�@j]�q�qDzHr��M^��w��B��⏞�����Z�䑴��-Q��J^~���i�/�V�����Ԇyd]��X�-�,:l�)uK#�Z�c?�G~>�-��R�@��t-��a�Z�_I�}Pa,k��n��E���$j�\����uD#+$�
7>�],��<w�� �X }6�d(�s�6q���G/�#j��O�!�G��w����E���
h0���8"�S{$�-[p;]��@���sQ��<��y>D*:���o�8�SxmO��V�O�$/3,FA�so�ђ[ �ir��/7��l����p�H�l{��zZ\��]A~�!|�	v��ޛ��_���5|H���j��$���o�s���%�a{��¾�����q�=A�J/���Ę�v{ ���I�|���ʮ���M0��I5M����	�I�N���~6"e�!!��rH�5�p�1��o�(��!x6Zp�����C���ۦ���i�sA)��,2��LϦ���a�������2t,?ݼ���rW/+�.�M,$�R��K�8#%��������$C� �r_�-�a����ռ���"FZts��j�EF��F�Z�f��܎?Z��hfo�D��_����!������`1��*?"�-��N�9���b�T�Tƥ��^�����	}�$������o��*�����'�:z�Wal�X� ��bE:�"�\���5h���������4"�Y��
�ÿ�L����V�ȝ#�^�>�d�/�LE�C��$^ی]Ow_��ߐ7=�*��#�d�������;���u�[�`��1ԮSb"r�ْ)�7����{N_���0��P)a�����?a,���-�$�r�\�z1�Z�7+�¹5�İ�K�t�1/�56������}�46�#����%eqH�����W��%��7���ōx�:�Q�@��$���I%�����Mu�
g�LdH��#�T��Ю��%1�ܧ7��h,)F�?���-�@��$���N'f=�Y����r}ͻ�;�9�.��<Np"��a����^t���Ϟ��P������T�ĚnuFc��5���{Ѹɉ�2Z��l�x��eA嗕9�
vE`+ggH �S��%������@K��҂�3��Z��6�q�)���5m���ax��e�Y�Z_�4��l��㳬�E�齈gD��r��c��Q��+doף�Ex��j};!Xىqb�\�}&�#�v4��N�n~S�&�0�|hA�錶�v��V�[c(ng"�ܮwwA�p.)�w�	�b�T� /yYU4���8K񃃺��_~7�����2
M�Ėd� =�/�6/)�&ԥ9�����U,iK���t8 d����M+<�l�V񄗮���$.,��(���+S85��˟Ҫ�6y�;� Ad��M�e��iޒ���.f怞�jlq���r|\�]O���6;*����UD����_�$fr���W��C�X�����$��Z��B"��FA��]�E?p&u� �Kw�J�����h�a�_��܃g�X`:�%�> ���q�[R��6V�D�6��s\�X~��DFhinI5Ȑ])9L4C7���y4���Run���?�G��I6l ��­� ֟����VREgbs�B�p��e3T�L��rHͩk=��z�tĉ~������Q�M;�^j�f-�#��l�{��ȶm��ِ]�̜�aj���7����~��}d�$��e!�@�$�f;�,�i.��]�
f�[���ǧo����7��D���ͽ�2^�r��R����|�ܕ��^���O�F��~������A�X�G�-��pn޴R�i���~)I+�h�h��B˙�A��/�=�$R˕�}Sd�m�-�Bc]Џ�����nbAY���������E�'�nJ��i35��L�k� �
 ,��+�wZ;�Sm����m��N��Eϻ����X3&��'�o��!��$�GǄ*i��?�}Ow������lh�R�{�LMYE����F�6�T���K ����3:�s�u����`?���u9s��E dɕE�zVڐ�)��H�=#Ԃ���<ۇK�b��J���?H�y�sm��HJ��у��݅"[��}����]�Fs㊫p�n�Rh7pڿv�k�C�ݫ?����5p�P� H��k��?B-��9��G�Z4C)m��:��k��u���f]H,a�t�R�"P?�'�9Q%s�"��F�l�d?V��<�b��(�a$�ct�-�
����;��^�[�:���>d�:�� ��V{*[I++�_&��J�G�m3����1?ˠ�[����7VI���p����ɳ!��Ć��X
��v'(߷�@%N��T�9*��G\gBx�
�M�	���p�p��V�eJ��N�گ�YV�G�j�VT�n^RS�%#sy)��Y�瞻�I�<�]}�"�g|:&� �?<������F�;�&�p���W�oY MH8��O������w�v{�~h�(Gg2x�4|���=2�c|3h#�-� l�ˡ�W���vg���R�55��.�'j��)������p�V]$��^s�r�aeO.�u���`+12��P���K잿�(��=�g����8����=��F�A��J���N�WE=���� �d��wu
�)T�%M�-+�V-S��J�a+(`ͧ�B���QMUX�9Liw�֢f>�h�Q�ʜ��fm{�;ZőL4ʎ�=pe�ߌ�6@�v�=�Yޘ�!Я\����:���P�J��r�	u����qGq .��ѬU����	���"Q<�iơ��Ь�@1t��^�o/�e�~|���\Ä �:���/����%C�v�^K�:q�"l�!$��e�
^8�<C���wg�,�����eY����-�M�\�`��ѷ2��կ�UF�B����v%�r�<�-��,��p'�"��Ia~dB��=x�qf��\�b�!�0�s�	L:�'ֽz�KC�DbY6��Xh�xl�Lz���u_�<fhL͈{g����VZ-�RJ��d�/�	�a��S��RH�.�-�(�UU���Vіw�l�w�8I�,�k@u�{bO��b��.�pp���9����b�����RX� ;yH����y��O6�\��nH��3�0b�%랖�is�K�Kb�:p�Z���ȹfi+�*@�#��S����o�����+e�.�_]�O�f��U��NZj�I��v��w�t����� a�%���z�����q7�އ�:���=,�'`/%�VRN>2���k� Ӓj�U�E�r�E#��U��3+@t�� o�yS�
����Fd���\y�ْ�bgroe�29��y���B�C���¯&@MN�����S����8-�C������T-#חGj��ՙ����%���mqvqS���Gt�,Xj�\�J;m�u �''s0~6y���g�ĸK��p+͡v��U��%�DXlxV65EB    2dfa     810�������eE� i�ݶލbH҃� �k��M ��m�VW��x(N;x�0�BK���q�Z�����+��I����A�[:�^�����F���*�HƢMO2��y?��ӳg��tU��� ���C�7���q���DO�����o_?��R#f���{� E�BERH�\��^u��^%�,�TI��V��{���	ս
��53(�-��h'G�[�)����Qz�d��$���8�/�����s�����]�\��@DMKBy�`����Fp���s�pDEj_�Zhy�Q�_y��=bfa��b�?6,���B_HA�U�:�^��/K�xl����P�6i�2b*��c��S�uFH�z�n������DJ^�U�3�Nm�Em��y��L�kS����6�Jw���C�^0IY��B/q�N��zI����w+q���cx�o-*��mm	�
3��I�T�K`�͇8�7k�5�ĈgnD多JG��g�; (D�{q�u+��k��[a!�Y}�a+dU ����t�+�Z�X��5q��zY�eb*h/o�r�0;MC��_�$f�Nv�H6*�1n�Lf++T�����7����;%��c�1��7��!J�|�f�f��r�����2�k��`�n^��_�N�j���p',BQ����E<�,�)B�\�������y��^\B�����R������;����1K�$'�]ٿ��A��+�U�k"�>��bFA*uGT�8e�)�dx���.d}G�<R'H���O;UGr�C�M�S²�k�4�T� ����?��Wc��Q{V���r��<�D�f��)Rw�������D��xn���G��*����E�������	%��{����f�	 ��-��,> ���>s��t�Ƨ*�܇����<业M,_F ��Mg~�T{w��~x�mV�o�aN�
9�\O�).� ��D�����FW`��`*�#&�Z* $H���w�g�(mz��3���_� �:½��`���א�w�D^?#GM��8�\��cWP��yP���~0�UD�����ݧ*�s�@��;����R�ߢIV���+����B:���8j�ɻ�r�yP3���75����v�
�4il��K�6\Č� w׽�"��/=�^L�YB��0�E��3l��d�<�_Z��j��;H�M��s'_���>��B�lF7����}����t�ݲ�@^N�+��Tp�}��,$!��o��������6���c����kO��oo3�CQz����#+ ���oߟ�q�﨡���U˿��^�H1W�g�]��_X
Ɏ�yK�r|�z)w�l�R'I�����
�0�"�`��GnO��8C/�ң{�3)�'Yi�{6?q����c.|�U�r)ƜD/D&��U�\��,0=�Y�DD�����gV�H�U�$"���X�^t��u�^c���Y���|��Dn�����]N/�|@v<,6���Jr�SC���D��<�G�:³d��
��#f)�@�
r�t>km��QN�_��d�Qm��Z��n�n�'E�_,���AϿ
�݌� �NBة�~l����<���O�F�[�l�$�9��#+�����$����.���q�Ƣ��h1�?���(�S)6G�v�Ni|��T`˃���a��:պOC�qc�d��O1 �1��I_&B�)��爆w%����U�,��.i�	ά��`��d�T�PJ��� ���
X�2z�����E���ϸf�Zߥ��v֚��L��x  �]�zU�E��\��%�b�K�pV�G��A�
QԜ,�/�*V|3���.0�6h�>N�.�+�P�-��g�~���=T�&��ꥀ0�n��o�3�6n:����j��6�D�=0��Ѧ�����i�J�'>���hǩ�t��u��I>VZo�	2�7��xEQ��"�e�[ ��}��8��~\;����3���=�*Mď��?Ƅ��V�(��;�fL"KW~ֹ��q�X��Fz���8���39�"�I*�ٽRiV��
XlxV65EB    dc61    2950�� F���]S�5�n����8��:$���P�~CBy�l�(�FD'=�b�����fkRnR�X�r�:���?�x�E�^[C�3����[��	6� �'�B^��f��j�y1z�{��V�t�A��S!g�-�e��� Z#�"�?��p[��+m?om��!��T&��ar��o�f�:�6h;�8�^'Kw�ߓ�y'��Ű�*C���j��l_{qW�E cy$�ם5-�KR5�x\F�����.46�Ub��a�⻍5,�>#��*z��w�b����{��ǝ�����P�2K�+&����X�Q�X�< �k��"��h��\@�M���K���aD��8��[2���X�ʈ�(��y�DD��^�* ?��Y4ĐP�7�0M+Y�!�I��~��r8��S��1q�����9�����,p�\�|��r��F��:����\������MY&�zD;�t(w�NQ	�-޾
[����)��.:h���O�go�j-���G��N�`�+����$i(��:�)a�貧C�\�G�n]<C�}��K��H�bq#����?��4n�oپ�ة�y�.����`�V��cf�*"�2�`�e_��;Uٖ�!�Oə�$��Y^��n7�F}���Oݸ�a�)��[Zy:�&m�Mtn.�cv�E�Vc��^!x��M[a����j��ngi��Ӑ$]�CgD��d��Um�D�1<z���π���\� ��y����&�xչ�5Û8BR��;��~�.hn�?�ֺ�9��\��T�k�?�0"�0�߸/�lAƏ�@/?�:]Ale��Rw�_P��g���_R�:� \`�e)�o������f�D��s��^�C�v)(� cU�ez�~�W�!MAd���Zm,?�6���Hu�������W��T��E��M(2nvi}+��ub��`O/$�VqϸtF�F?%�����������A�4�]@#uu�0^3)̭�'�/���+�U���s�<���zp�*�{$���#i9bF�׹�ʀ�c뎾=��n��l8�~(�/y����f?�	0����~�f�	Ѕ��}�Wp��5�mf�NI�#i���	œ�7���[�����`<�n�v+�Rm<��Q�U��ƪ(C�p�Hʪ��^�뫁�:�3�$@�0��l��ȭ(�^�N����&��$E��w0F ���S��n�h �8���+)��y�S]�tgߧ$� �O �G0%��O�#ņ���������?i��b�<7ڶ�{j�E�C� ��7kuW��A��B�#b��W!�������C[��f��3y�J}.=PC��I��nk�(?��i�1�4���k�#��)�*�����A>��  N��2Y���6B?9����dn)��z� #h����K7�u�!��Q?Z��~~���Gb;���aD�@�Łbvk�	����7�+?SL�.��Ύ�?w�Àà���H���#�Q�@ć5��S#�O��� Ѭ�/�~o�e���QՌ�~�#��0���'�d]Gi/�U+�p��/��%D� N<s���܈*=^��%��W<̡h����l�.�uW�WD{j�ć�*m�:e�Hf�Ԭ!��L������(���-HG�}چq�e�a��\�$�oV#�$��Q$@����%`V���A�ae*�������|�����[�o>Ij@j��j'ñ�#�����=�k�q��RA�0)�/nbX��Ą�0��r��B�����)+a�>�3�Uz?�����ne�6�E�D���|�ܰ��p]�F��%���0��
��R˱@�Ʒ��}��P��k�\͗����ӡ��,�r�)��P[r7ߵw�8�E��?dR��[\j����.�[��RR(��|L�WjZ��o���-+����u �d�)��6+�kcy�<F?df;�1�Љlv��z$BlKm�TI�:D9cؗ<+�����6k��&`GR�(��v�U]��Z��f0P�^��T5U6C�Q�H�N�&;��쉹��[��]�/��͖����e� (�w�K����{�B��(FA�Q��5���M��ogT'$.-���-^�i�j0�
�	Ӵ�{8=�pe#�@AK=�1�[���")E��p�S�́��Tǋ�������:]��g~̻�Xù����ͱ��Y�&�.��֠1�ntdү���&LO��WJ��>�b�d8�MQ~j�X��6p�J�</,8/O@G�<�������s�"a ��Hi��/Am�,W@�Ev������Z�u���%%G&��E�,z����2S9O�E�[��9�@d�R{�Vu�hL��ǭ|�%��cS��kY�)C���X~��Nѯ>�p��=W�.bjWҬ$x1�Ʈy�� oN�
['���T�cS���
�E��H���̄��s���Mt�<�PLZm���w��0�/O��') cR��Ⱦ�2⟉�$�=  =Mee�J�X�o_W	A
��/!�D����m�!`k8����Vn73�\Z$z4����D�s��~�E����{~��]̿1�k��V�,�l$t��+T~mZ�_/g)��B���"͛����Дj&L9�H��L���#£�I���{�n|�ʑ.�q?�u�/�z��r���A+@N��M�s��K헠�g*�kn����=�=`����G~Ԇ���(�ֶc#��vg�<)�?[�ci��XaZV�\�4��@jWb�pF����:��� ���u�d ���l��D���jq!���/Z�[�����g
��n��9�2P&��\����T]y8+@T���ީ�k��L�ժ�P� yǮ#-fX����*��s>��@'t �)��d��X;ti����D�/�s@U���u����Q���Ӎ$m= �d�I�q��T9&ɖ��ѕ�&a�!�?�lx�Cf��:���Nc�~�fo�:��C�^Τ�	WH���1��A;�2��t�1��G�9���b�����I�-Y��J����#kc��N2ア[�L�z��ћ��c9ز�l�����7�S� 46f�F��!����Hh�۫^�a�n��5�и�~n�7�m6D��D�Q���K뫄x�[b�"޺ny>������u�~Y���M�4�HM'vM�&u�4`P���o/�ES�C�C�ve$�%���.zq�JSߖM�kd�v�4�+�}Sc{�+��6YF=o���!բ[d�W��+3��ftAf��>�v��G�W$�**Sܑ)���t��X�ܮ�#q`ZY��颽Z����7�)� ��Rk�m�s�t�$����,�;O�HV9ɀ�E'\8�9g@]TS]"2RWAx�nN�m��A�H�����C�L7��o��9�	�Ԅ��cɂ� ud�_j2/)l�m�p�(vg��y��V��/�A9�wN���?�Q߿��U	�:^iU
H��}�,>/ =��rx�q �k"Aû*���:{?��&�GW��I�ͳ*�E$%uy��Մ�Q��c������������~�5��
'�Er<��AV����Rɛ	�k������W[�N�'���Jz?N��6�e��1hcp3QfiR0t�ư��|.C��l��C��"���9�7� �=��X�n�fQ�]��T�u���L S�Q�K!u���q��)�ݐ/L�q�������p��1\k��n}�غ���$\ê��7
0w-g�ZGP�,�(ʘY^+��x���a��:�E��D��u�(gD���dF�Or�U�+|���E*����j�T6��`����MX�3��?R�V�o���%�*��;Ղv5K�����ƛ���'=�RL�y��I0#N@�/$r�M�}zz�R� ���a�00޺D�w΅�ʀ����.K�G��z	k{/���J�i7���x��y!�拴q;'��Ϸ�{����t�������yƼ�@�굀r^�`G�0<=#�W��}�E�>Vt�y�_>��V�����=���O%���$�G�{+���&�k�����b�k~�![�݊��ΞpE`{ �;��x��{�e#�u�����E>'�Z�7;�\�A&7x 9|�n���h�؍���K��;�	�����O�� �p_�2;F����C�_Qˉ�3��w��@Ƭ�~R��L��5m��GV�"kFh����1�PjHH�;����r�a�^��.ޡ�ѭR-Y�A�qE���͵��
��ٍD_L��Lы	�n���&�4�_��x�-x'{D�9�<d��أb������ǎ�P�'���d UA/��$OD��u|�5(}+y��.ʀ����I7'5�G�z`2 �5���`H7�C&��d���8���3re���:�)J�'��4_�v��a��� s�NH\1�L*�}�\��A��]�U@��d��N�kf����p���,Z�~����K�ُ,���Z�WЁs��Z�fU6��$�ԝ�v��fs���	'o�7
�Mua�AN�3��qH�_%�H����_���MD
0��u�jr�4)����-�K�T���R�z3�p����A<(@A��iz0 ��w��?���W�_V���b�PX}wLpMQ)͡A?��k[�m�a���M�䗋W��,hDѱ�m�9�0���H.2��t�v藲L��ǟ6�DKk����sh����>�8S�6D8'?|$A�n@��T�Lw8��+Q,���fp'��9�������H����#��$��o��~����L�Y���$��w��=��p ��J� �׶���ttIt�"�Z4�:��[b�VΞ{��}�~��) 8��"�-��+��9K;*�$��i�}�!�n5X܏HJp���L��8;�s+ɣ
�_9�%ؔ��QJ��P������/�	�(���:�y!�����BAc�*e+'���T[<gw�v�v1Qȡ Q,�R������,��1�����B	�t�����T��@nt+�WgA��o�1s��jXr6����#��N/����݆�n�����t5����nE���3w�1/Wrٷ�}cǆ�Z]�I�v���gI�y�a�\x�2�T�&�A�`�ޝ�Ҕʗ�ީ�x(*�&�k��!�*�nKl�{G��rF�Kr�%3�GL,���	3p��Ā�2eYΡ���5��!Ϣ`$|)��� �-��W
1���e�@o2ⲴRߺH������t=��=�<�h�1�~}��	�򻠷�.J�q��������MQ>U���གྷ�8đ��4/s"!�R��/�?��G�}^�^�ތ�����f��z�,�}�%C��e��������;?%�ѥ��6��r�"��6Xϛ�NIJ���2Cxs*�cy]I�G_�G�2pܹ���QW�AB����N[n¯�u�vvH���حtX��*��
����9���۱��Q���=�T�_g+�?>^�j�6!Q�2�2���0�l��ʼ�"my���Um�Ai�&负���z�e��'�X�������T�ʺ�|͕��nx���W�%��mǔ+{��E�gL�2ul�F�4y��#Hׁ#�����]4��h�y�NX�zPq}t�� k{�;W�Z�"I}f����]����h]]C�#��)����O��V����9
"}�	=�_�je�6Ȑ��u|�~"�љ���h$��2uT�ip���b�-�hJB\[[ �kij#��
"c&��/��)H^á0��賃؄ M�]��':�ܔ�5dV2�CtK���]A7�u*��eLK�eiz������<B�Ņ��ۈ����@q�P�R�_3��m�ٻ1��s��m�,P�y10��Cvaj�4����l�X)����F͠��,
�u�E*�����N-�7^�V�rC�\���Op!��Im�� �Ve�����X�G,��߼�A��]��wxm �"mݓ��%���KH�fdP,�
���E�yl�u,9�v�M�7�B���'��gIE�bPw��*�h����%��l@�<�����e#�Zc�T%�`#�U�d�,��37�\��aPSB�k��m�
i�����^0A��'���]���A���H�yυHI�j��w���G��`��;l�N�3p�4��C��`��~l*�JNԿH]��?�Cr "��ͱ6k���l0��⛌5����sz���/5�(�pOQ����&�6
%�դ�����	p���IC}G�с�c�X�X ��L�)y�A0�E�oA�"�ce��l�,
�AY�����*.ELcu����ZͭZ��U�{�Kӿ�_aÈ�<^�k�C�N��i����k=S܋dG湃u��/�����=(��>#���krJ���ģ)����L\�,��b9j0*$���z�4�
��X4in�̳����Lw��H��B�Y�zW��̋�1�$:���|�>�N@��V��1��%鑱�| ��2=��2A�uc���.e:�AcTG�a��٦
jН'C�9~�O�+���"�D�ca��DiV�P2�M-�E�ށ'Ӵ�� 	x퉧�����J����t��׬HCQ��,����@E{��v[x]/��6�>���%n���#�l�݌�b�T���&��B�ě
�ZN�l�2�z6̘��;�sF ��
���g��}Ykr}�>5m1�|�(��.�Z"n���M_� ����Р]Ѥ�yY6���r���$�q�@/�^� � �ew��»�+[���@�G�o�a~e��oL`��a�_4��q��V��4�g�@��|��m;��@R'�\EeF�o"0b�"3���L�H����F�b&[e�sN E~���!|AX�A��'k��R]�=���M�*��6��Z����<��qL�_�X�5E�+|q�f�.ЭN&k����a��Y44�i����\���������=N�8rP��K��ծ25-pfN�Ed΍ԽO7J`<�;������mGL��V�7��9���ӎ�R����G,���R5
T/��*�,�p�KiF�����'�ӏ�2��$(�KS��9���3�x����M/��eb��'���u3�x*�ʝ�#�h���ǋJ��G�O��q�-A�a,��/Id��/{/	E#�h' �n���=�P��(��z�c��mvF��	?�7_`�S��ƅ���I�w�O����*U�#�r�Eԋm�����$ba��l3�[�������}�}1ѯ�/\y��1!{�iXR?wF��Jt�"B�fJ
_bf���.�����ӌ.M�����*�P��F"d`�^��+4ɞo-��(���)i���3Z��YWikA���?�c%�<�� J�k�g�+��T�<j��j嬠b�<<hC1Q����3�Ƶ������ ���i1����ϰd�F�}-�m_�U"�q����ڰ�F�p��PU6#ȃR���g� ����>���ڇ�{�e"\�
������-��ڈ�pU��h��uK��}���E`eA��BS��5��ƴbȓ����-���ǡ�)b�v�>\p���w�P��]�a���Ffe�z���2�����F1����R'vח�Y2S��'��c�8�b\$���Q����F�8���7����b���8�X�J�b�!�j+w��R�9�@0���6��Dg�ۅX @��_.��Vo&)w�|��W8s� '���fRu �ra�d�4�c(�����A��Ds���*�>F�GB���p��_ ���U������$<��vp�=� �U�u�N�a�c�@�[#��ǔ�K�g�����(�u.������u�o�2�b!ә�׎Iﰰ�Fa��%�*��5�kk�2j�[�?L�V��M~��vy:ub%4��}&��ɩ�c�n.�⬛�	`�����䫄d�^8���vX5z+��z��}pv�<�JS���_Kp`HVۚܿ\�KT����D�,�ئN9;��P ����mF ����c��+H}��Np���b�$���OVΜ���q��i��L��B,�<�)��K��e���JE����f�7k�*X��h+E��
�!P�A+V�!T[��y�r�UZ"�l�r�f�u�1��O���#��$RU�ށ��@7R�v«?��Ӛ��ũ�X�$S�)�䝔���~jns;���P��Q6����_��TЌYlF �DHW���"�@��oۻHg�6\� ��:*���#�O�"�"h��fR �����1LQ��h|@܎��6�T���)�a��ꂀ�
���óޓ�%�E�����*t� pg��l���o"��*M�|��\�aMq�D�׿@����ۈOW��l� [��YܻeuU�����E�7h��M�E}�7
�e�����$W�[�7c!�i��I9������1֋�w���.���9^�_=��6c3���QE��QNf4�{Mv��"|fM�+��Я!or�0��|B'ՠ;���T�x��̶� �b����V��"B�c5�u'�7:���6D��[`�=�D��
���m�WpMY����s��"6V��?o]g�/@�<9d,k���qǻm��q	
�V��g��P�1���$���0�����Ct�O	�~`�x��)���hy�SfE�8�#4<6֎/ ������E}T�,&7���l�bO�|K�+����"O�:j�����K�m腫#�Z��I�9�I�G�E),�=��� �^�PG��,ae(Ҕg�sj��o��)�ѯ����~g��ä�a��V�T�L䘰L�O�T�*�Wz��7,��v4�]0E� @�
�C��W-��6}y%���%�Dz�N�	�^1Ɔ.
���>�ź��]�%�'2P^�^V��?z;�� 1]T�Q�����Sq�k�G�e��ȇP���a��c����R�,����=��aDv��� Y��c�F�?���[p�1$���jC�|����0_�]����8��-r��	��]g�����: g��gM W�5Qjt���狿��=��}[|�E�U�	�P�̻|�K���G,lY�����=5q|���c�~&���	ǜ4���N����DsRH�Ay3���������\���
%!�z�`kJ&k$�m��B��U;���t�`�~ 4ی����Q�ӷ��0m��@��)�/X��	����YT�R�hd�{*!���x�kf|tJ!zHB1�E��9s��Q��w�s���/JUj��y�]`�29��S�vH�ڬs����5`�8�#�7�e�>>/����Ÿ~�hi�,i�k��x���x$45�C�ơ^�ײ ���\��9�>o��N)�x�/^Wk�εU�Y��ח��6��Y�����w���.�	��p1myq����������Rk����i����Y"��G�����~}w�7���F~��H�@����~�����v"�J�*�����	�c�*750�0�����H�C�G-��/cIV�0:
�9���{�����Kq}�v
�z�-,5��+S�!��%κ�ƑlF�0��3I�c�����B�� 4{EA�aBC��}���$Ѫ���}���_2�7�}�(o�F���>��9���~�;����-��\G�!G)"H��~�o{Ȭo��т��Dw��]���5+�TFZ]�aG7+�GF�`��������.�9r�qX������
��_��׽��#�9��A�b�*� \�m��Fs;�P�6P4��Y��7Z|��0���I�)�/f�d�����id�	@&2�xJ�;?�d$�T�P��k��:P=�$��=���#��/��0�F��T�:i�%�h]�K�|k| �*T���!!䤌t��/��9̖�s�jd�����F����XG��W�3P��ME49>9�{7�^7�+��+��g଍�.7{��dc�7�WX��7�Fh\"I�V7��1��qځ�|��͂�����5���h�^���K�9�ؤm�d��j�O~[Xж�<�=�'&#|UM����]�G��% |�2� �.-��������c.;B,�{a���k|��D����y�	cY�gQ�Ĉ��i�b�4�BI�8�zA
w�*��0�L�]��{I������4�*�U���X�UJ黙���s�ĝ�]+���0Q:�.5�_�0�/"%�s�dm�@�(��^A���B����*>5�ѧ��dP�6�[6GQo��A�MRY�q�J�زUɵ3cr����s�;�������Yc�D��ʓ5ض�lVɔ����.s�����e@�}:�ڨ/���`G�D�����	s�Np�8�d�)ԑ�)���T�r�\���n�g�}\>�7�1^M6.�v�bV(|D��@�8}A��1+���{i6w	��D/��(	p�,V���Nk���V&{�)�L�c��I�0�[A�������Tw9-Qn��@
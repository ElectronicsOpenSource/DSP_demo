XlxV65EB    8a3c    1800y�p�.hS�8v�{e<e��F<�p�T�]DҎ`ɸf		I=�+w��K��ʘέ���	�gV>�B�KZmX· ���ZlL/�vzi�̢��+z�@��A���@��Pkye�ӱ\3&Z7RN|�6�U|�0�,�,�3���·2ͦ��-P+�������ڴ5=b
�b���uN��j�E�X��m/��(%JE���-�O�z�����q#�hn6��t��J%��j�_T�7'}��X�Մy"��:���9:�j�I�q�N�]f���E�g?A�ܼ	p&���-�E��9�qL�[�cp��3Ո?ԼhJ�&�W-�E���S���H�Rk��8���M��O�(�Z?*�$wr1�<�-�S�hom�pX����ּ�쇤���>�)GnYM��B���� ��6��.���c�
$��7z(��&ݏ�DM���2Oj���\�h�W5A9>�$�<@��gK�(v��=��S_9U-4%L;�t��!�]��eJ&�1V5�v�����_IA��!�m��p�ac����v#G��*f%g+=��4ON�u�'e�ӷF�x0e�(���l�np+8��v�/�5�X�w	�ϥU���<��va����P6��Ԧ��x���1`!����K�s��D��fZ=Ǥ��d���t�q!{2\�"�>n��'ze�pE*Ŗ��7���{<(�L���y[y��;1�d�IE��ɯz��R�m�w�	�B�'3Z��p�9==�>@�E�k`��h�K�����Ƅ!�:~�(~�d��g���7ac�?s��N<�Z��@��8Vd�u��]�7�/ب̟��N�{]	�˹�6 Q��17��y*�Մ�DZϠ�W��FhȈG�զ.[�{��U;�E��=���T�����G�(T���CǇ��̛#�b��#Sj>Vr<ؼ������F�8��۲+����%We���V�cO���]��a�-����.����TP܋:XlI%��|)�t�<���٤�J��8:6�9��0k4�]��w-�4�f)��$�m�Q��J�B̍л�༮�e�{ڵ����'����\�	��+���WY''���3\P��6��>
M��X�L����]��E'���� �c�/����5�ǝ� Uf�S)����}=�-������5�٪����F����
M9�[/"����9�\2@��z�~�7Pi�֏�B0����#�v��Lg����X+(.Ք�cZK���������y*=g����$�{.�b�E2��ub߮��?T�� ll>�Z����+e�Gf,���T�T�D;îX�<ղ�&+L��e�]P]�����yl
'9�XnY�ԟǘ�Kd���'��Ӝ��5�#�׵c� ~� �j3�5�==���+g�r�
T%�\?�y�X��L>	�Ցk�)���d(6�G(����d���@<<`n���Gvi��������rᕢL+Ô)�d.��q��"��Ɨ��rH��K6�߰i����'��G5j��P���[	��ʋ{(�<�x��6�sq�,G��6v��ڦڞ]��G��<�T2��k2il��
E@ �g��ep���`�!AX$�w:)W��v���P�%�L�U�/��p��%�nr3?��f࿜A�f�����y���+ꇦEŜ�[����IsQKu,y���6�V����&��/~8m�����'�ʧ�)��Ţ�&���ʘ�z��ڐV���?P~0��\\� �B�J���rvn�	W�������hY-���ÖT;��7�Nj���Ǭ=�O90��1�����k'�qZJ��!�����	��w ����'�*3��s���9@*ߖV��@x\��ύ+"z�-�R�[��A�,�^Ӷ�qzp6��4��7ڂ�@��! �c������tP~�$�X��\\��J�HR� ��ێ����?w�Tl��Wdd�Y����+�O�@(!�Fp�t���I%��� Y�*%Vyt���L}���e�V���A���x��Q�9y��Fpc�u�!7��n>t�4���_ �7�ɟX�����
nU#������:��AY�S"��|�©��`ܩ��:<:d����.�#���
aXX�(Q%{"����p�@�={���r��r�\�j��+7��;遂XB�lzo�c���u�F�ie&H�-��q���(��%)�J�n�绀� �0hTڬ���BVuh��nM�@\�#�ס
�¯��`��O��B�p � �k��1���;];��u�C���<�;����G6�M���g�0���oL�-%(��-Ghn��K.)��/����OF�n�F|�?�)e��Ҕ�8+0�5%��|!`����������cԴ�fF1�d"6[�ܫ�G�>�����T��%���|y�ǿ��H�:M��'�ڊ��	�e�h5�/:뷅�����a�z0}Y�F}���;�y�J#ag��q�!kt�u� l�8-4w4��=C�x�52�D�'��4�@�W?��4=�9e��0�x�C-Ri\J�y~��m�_cH)��r�c�U��O(���%�r��A�;̬i����VZ;��Ņ�A}m��j�~���73P[�P&X��,������2y��Gm��s;��lF<���m�+,τmmO�����[e�3�n<"���A�@�[�};���	�D�ؘlӮ�r��J,�%���P��e�P�$ �mb;[�9p�����魼�\lט]���&�Tд�SǷ\#Dv" ��H"]��v��$�ǺԂ���cP����%��xǑ9�'O�.�P&�gK�N)/�T#Km!��|Y�"_[�r����7����;�fh�4�Yi�n��v;�~���1]��>�U{�v�Z�� DX)���w�̥DM�d���r�3nnM���+k��L� wK��J���1�	X��SM��;�N���)JG.~ˠ�2c5׻��g�/��s��d�8�@
@��\��e�}R�k���Х�N��|�=HL˜VW{�`g��-�"�HE�,O��H��\���wND�ilf�OG�4]47�c%�
ǔ�g�ihl��=W㟦$���V�����.�J�o+2��oV�񇯬���̈rB����Ψ� .� ��-����iK��y(�zm��qb|���iX���F,����'N�G>"#9@`�l9m���k�K�M$G�8>T�;Il����w��w��	�먘��l_�ng��S�H%�Q�sS�_nD��$���ԏ'�_�=���Dh�{m�_z�X�K���CQ@��hcסfRy�\Љ�G�5��M껍�7�8�Vޓ����)���ۻȵx��ٿ
�ˢ_��k�eO�A[�1Ӧ���*J��}Sj(>�w�q}�<s=�����1���l�!���V̄����������]L���C:�(�E�t��|��),����Nn�Pi]��Ll����r����_g|�D�Ɛr�r�#/�=� ,Ѫ@��K5���Z����5�O���K����"9�}ȯ�#�CI�TV�M�c�����k��e����Y4�evH$���(���� -��W֧��':�!LtcԎ�{$A{At�AH��-��/m�ɛ�E�}�56��������o
��b�ų�=l���v���.�h��-��0e:�* ���i��r�W���D���/-{e��C1%�a��y�cD�bE�����.����䚙R,r��<��@����_��aY뿊�o�[eB��d?pB�W��5���Q�~��/~�Ӵ	��?O=ք����م���!Z�R�p��6���J�t�6����zk��ϫ�.�H.����a����Ml�8�7�+��:�[$�J�_��J5����Hܤ��(S]�MV���p
ز� j:��j�@H����>{oZ��Q��a���ᢥc!���j͎¶�|}}��^i0/�����*"��m��$��-�|x��/I�N9^����@�Dз��yI!jL�T�k �)LJ!���f��fc����K�Ґ�dMg��U��MW-��:�����&�����%[���NRt��)��6(:��>,�&.��/z��ҳ�y�+/6�B�Jʳ���:�b�/�B�cH'�#�s�l\}g:i[�������i��Ϩ�AM�Ln<��S�����gѦ\f9�;��D
5=9Β?�!�c�3�6S�Ī�PlNb�����cz RC�СTw���?wC}��P�JĎ��i޹D�Y�`���=�<X�B��ɿ��p�2t��\H�(��v\I��v@1����_	Hw�x�P�z΅�	;�&�=�,4�7c�Bkg6�c	�6��|�qu����շ��I�[O�/�Xg:�,+�9v<7*I���=J^{W�<�]PY)0� �h�d�Ks[���_bܵj_���r��~n0��W+-�;~���"`���<F5GWO	�ti&ʐ��R))$#��9W�U��w�
F<��8��:��L�Cz&}�N~��hf٤���l��L>�Q��#�,��X�[�e&� �d%��	���#U~uy4��1��^�����TN�Ӆtfo��"D��s'�T�C��:�ۑ{A���������!Z�R�^'���f��z�BP��Ec�6��k;��"���ou��%����+��>�~��'�D>���S8���d�]��m�s=%�}S����!���������
 �zA���	�gii���l���rx��C0Ͱ�C EAiFm6���J,]��C�X�\O�Y��d|�Bet\(6�Z�=��}�R#���W�����H1��0K����.��ZȽ��j2��@2�K��'c�L6��x�6�*��ޥ�M�����Yd��L5�ɸr�J ��n��t�R/X�����O��rOkw�P�~+�I���^tr�PS�ޛ�]���hܛ��D��q�'~$W��%�#w��?z�a�L��ng�R�c��Y�b����������K�)���f�9U;�+(4j��L�\� ?vY@�o�{���[���q%�H��nj�Lv^'�;������~z/�ݹ*�\4�P���z9~�\M
+�h��HvO�����B?SY�#\���"�.��L�*<������+�#@����t3oLS7I�Nz�Ć�u7YXQ]��_��z��a��N����'>�yj�=�_��we#��IDJF���&UX�ґg�X/���v6�;�{�6�c�\�A����t���o�Qn�@��N7�<h<ɨoad�-P�?�q?�I��+�bhHf�#ӹ'|yp�	O�������b#��4�(�^C�-D�I YНuKy�;� ?{������a~�yK봟wu��J����k܂(�Z[�Ի�����b���~���}�P��!0e�K���	��P�R0Yy�6cgfk�=�[ l���;zN6&�2����'�Z�p:���l�Ϲ�W�[�T�r��)D���j}�ѐ�E��*��㚓�Ps�`�a�lK!�����7�j���5��<��V^���E��5YῪҨ'g��y	Ю�X�z�<�H[Z������PV�)ΌY<��Tv�(�� �sZq+T�_���Y�	���V�PH�s��?�7�4^Ǹ�� >hZ����hYl#�|
L����<�c���$� �QX �T�J0B8d���=%,*B��d����:���N�I�/jb7|!��ȕ�W��͗X���l�n���	k^gLoY^�2��jx���3@���6�`��x���{��MbM�������X������#�:U9G�j8���nEi?�w�}n���v��E��D��0kF�t��p�Z1۹4�d:��҇���H~2�7Ҟ�."�!���Ø�G~(Q�q�����Y��+�y��k;Oqs"r�,(>AEU�}G�'��(�O|M�ϙ�����`i�w�be�P"z�H���ᑯ&r #TgR�BR��2xP@��)4�ט���B��z���1}��f-�������U�N�ۇ?N�
XlxV65EB    2798     c00��P�ٙ'�8u�ozNDG�j���1CF�ҳ�Jw�c��(��(%\RnG`*���$���Y�7_Ȭ0j ��y)|x�ܗ�uk@y��O��u@�ިOx�sֵ���uq�$I%�Kr�޴U�{�?��h�C����^�sy
�<��؁�"��d�ᆏ�_�{4~6{�Ӧ?<;���62F^����F>��3ߩõG��G߇�Z������fb*�-
e�;)�qN{H�����Ü��	L*̮��,�����ʋÐ 
1�r��h[�ZP��8Cc*���<ш�	�_��y��F����9�����$���É�����!}�h3t ��R��Չ_��V�F^q5ō�*
�|��4j�B�M���Q%�3��xG���v6#���PHˢ_��m�

K����׆q��50`����������)�sV�VN�ef�)���m���F��?(�����s��ɯ:��c�B�V̮__#������v{�h�X��ҡ6��ч��=鉪o�p;���)
�x�%�r�8�KŏeUS���O��D����9hn_gl��/�����+�,�Y�=Rh7s�3�`P�R�D\��l�.%�4m�:�Pl#ѹI�:�4g�z.G�6�!���X���)��~{��%����MY��dT:�Q0����������$w]~MP;,>}�+Ŏm;!�qcqȆ����XRN�U�����̙�K޸
�c��W�'�	���ٷ�]/���ـL�u5�l^As�ɟn�M���a�
]\n�jG�2�:&Q_(4�X��2��Z���w��#q���P�M춲�����bо-5Z��Y�.��9��dl&���E~֫l�[�G��Q��w�zm[���l�[����`�WY��W��uH�͙g�}�H(}W��Y����8��t���u��i�� ���nW5^A�p@�5Ӭ�Ͳؚ���$-�B������K�=7���	`�d�2�M�j�bi�jSdKv��<نU�Bױ�1���p��o�.nl�d�D���7��rc���#nÙ��5�D�y����I��<(�H � H�x�?��iNK�^���L�+c��'��^�΀tp���(^ie9���z���?@�U/5����sRa_��ŵ��7�M����;��U��Ip5fR�%!����Z�ž}d��P�V��<��'#Y��5�X��<�G����T�5�޾�h=�;Ka+�H�;"r�bS<�Z��]���P�M1�0�
�W���z��7�jמ���4)���=��M�ȷ�ϋ���Ut���@L֮g��ޒ��g{�*9�db�lV��M.1�y�:%� .��3]�]I������s���}�"�K*�q+�"���3����(�
ϙ�e�
}|�`�=��Zqi��M�jt�P��t;9]JS�Fױ�4�������S �0��?�8�g��<b�þ� �������?*Y�i�Ѷ��W_T��U�����=��3��R�#��	�63�}ֵ�ɱ��#,�w��?V�`��Kd��S3E�ȗ�&�"*�>�(:ׁ����8�{iUn�oB��8�T�ؖ��pA�D�͗�˭%��)7M�tr��R��{���J��B��ɎB��9$��F��k{�p�W �9,����pZY�M�Z+��.�3$�yff*�~�]�x<S����
�8U�h�q~�4{-�P74ܯe檀 ����K��$ߗو��U�����C%�7��X���$�����6��uQB�%���#��	��Ȫ��l\e=1��;1T��:Gi)B\jY���"t�^9�R����E�f�.��=��sv鐏��ͺ6g������	&��q��O�q4�����w�4����L��"�{E(��/v���n���V�C�����M˺�	+��*�1WS��d}X��Q)8�����eo�r��iI���	r�)�j�� ���j����f������f�%ȡP��{?����e�5~�8n�[{���)�Y�༯IuӢ�P�\<!��b�|�Y��9�|X�(i�җ��SZm��ϟ?��mJ)r��4b�Gh^�A�����,A
aR�UR�ݴP�xH	E�Pb�X�q���KO90/�ᩫ?�
��� Df�8�8s"�3I�9V��Ǡ��h�Pg��o���H&��^n���a		g3��_�\�
h �i����2)�R.!� ҺH�j��qFYf6�� �Qp$#�q�y's�$�"k������?�D�|:{�g�hR,�� ׾\h�a㺏������a�2�����S���ΫM���x�+��6U:#���u(c�$ޏ�3���:#)�֓��K.�åR��8j�|���/?ry�G�;����[36c���K�QI��Јc���G��������1A%�c·��77F
Z���RD��>��T@�ם��Ԩ����:lͩ~R�mZ�Js !�������w(\T��!_�F#I�v�;��-y)P�.ϰ���+���۟��=Vk��
��a�A� sƁSf��T�A
�h��%-Q�c`�����Η����g�d�I�U
��?����Ha�@��:���:+����$C3iy�v&y*��?DM�@�={�֛�-������LN�����!���s��zĂ �/��2A.�1���$��� ��쏌�A�ʓ}�w���j\D�ӲȳY1P� ��Z�b��X��Ϯ=9����e�I��T��}����-��͙�ciV�wQw+���n�)	ﭸP>1f�#l7����ߋ��m��D�.�:�a��0 ���D��A��D�^��w[������1_�[�c��I�'�]��UI��Z[�4���q�f�
:T`cOA�+}����p��n9�ג�+՟Nkߡd��$k�@�J���;��M+��ĩ9f:z�/	u�:�oVy��H��::Wr*��@Q�ʼ>l�}����}k����p�{����J�je�'����"�Z��+����[
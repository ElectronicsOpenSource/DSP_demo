XlxV65EB    4fd8     9f0�
hv���AN׀��':������<a��L�m�T;�O�#e�&dG/��� ����*��!_�����w�8[}��d�������҇Aq�
�i�YyR��iZVb�Y�w)��[�����3-;��-�&R*t�t�����Z(��~����s|����8��N�u,_|,K�4��`	�23��PpBz��W�1��A���CY��ln���`.� w3މ;�G��G��cF�t�Zi�d�&�����Q���D$�7�@�}��꟏)El�V9\�v1J�s���L������}� ��"H���v�`Bng٩֏����t~� �s�ۊ0!M7P�<Pʚ )���M�>J��C�[VP{��k���ě�fn	��H���'`��zߡ��kjO��h�ȓs��R�\˪Ƿ]mu;e�/���G����H�����}����t�F]�6;��q��1$�S-��T�����/�a�XS0Ԃ�FW3O���������U������F�u+�_6������&Z&$qB�Qs|d>g�՗5h*H��E;�\:G5S�=���YA}�E�7	���ܕ1��K�������f�p�gt�
})���z�"��˺\tVV��F��YM����[[�Kn��*F�ܯ��5u�:�|�#��߲ː������N殦�(Ѧ����'V�9YkI})T��"*W�Z�p��v�lik����	�7L�na�����@���a����A�)���8<f}=X0F��6��{�)-FR�����ӡ�0Av��4�ċvY;J
~�\hX;Cf!G�xN�v��en3,�`�8�*�5C���0.\k�7|=�H�QW�!�f`y���i����f�q6e[*���!�6�|���c_�U�J����K(F>���w�v��y�khT��5��x��U秹 u"s�Bs�8�Io�^1�U�П~f
�e�*"[�ς���~�XM �#�-g�*g�>X-��F�Oa��`�F%)2gL��o`٢��=Q2�B�#��Mo�!{1Z٬Cq�C�
�5�*=��,Y�2�{"�z��5�nBR(FǨ
ѷys�E�$}�*x��R�����r���լwAX�;>�-x��f_��^Ko��VP�ٱ��.2и��w�I��/@��o��\���j�c�D�����׮}e��7�X女��,Qy�dǀ��� X� ���i��d���!q�������gG�~k�h2v�֍�9(zQ�N^ȕ*�$Jڀ�a�~zrV$�S�)b��%&�Z;:�qԋ��2S��L�v�2�#]�%Ă�1��A�
d�G{Kc�3����@�/�W&�'*�z���-���lJl5��ä8 �=".w�>�t�K�	`�%!����)\<��<?���L���y	C�-# ��pY�s�~�GS1���J�`�������i;2�-�l2�M����2,�-��+=��:��	C�o���Z����[��ٻ�,4#�
!`h��5{�R᮶e6:����4�Xn��-"�!
����=F"�z�C��O�؃��
ګ'�쭝�=r)��ʭI`̿s�-~7��Ɯ�]���[9Ƴ$�e��w�a��4��yE$��n��Ɖ&D��%�^K��e}�����W��)�'*�A���B�mv
F`��1��4� �8��pK�AH�"1�'m�SoO����h�B���#�3�t'K�m���f�H8g��T���[{3yi�ԍ`>ňF��ø�P�Urc�tci_ʲ%~:����;�O����a=�X�g��)~-dO��XVވ���z;\dy�-�@���������.���ٿ����C���9�Ȑs���J�wKp�:��SA	��$ǀSQ:�6o Td(.,LW��0���s��1|k�|���{i;�ǡ@��I*%C���Χ�e	�W7��|LG~��U�!�����i��魳�5�#C9���　؟I��ʹ�׼���ϩ6�vyH��Z�/􈉆��ӗ^�{+k��^fҀ��5�D�I#8{��Ù~�9?���>t�n�@Iq�V��+�z���j��p����>Ap����e�����i���R��8y&�R�i��>�H��63��&��S�*#=��Z�3k�5X�Q�w�"՚oR�4�}#�a�W���<q��'2x��]#Qך�ZX��[���>�c�P�����Z�y�P ��	"�T�+w7�R4�9\E�\�Y@�4*�>�f���#�j:5��7h�g}6j�UX�T��Z�u��xIN��I?Ss�]7�N��Z$d8���1�S� �m
��J�Y�PXN�{�y�8���d�w11��L�7�
8���Q:fx�~�锛���u�Q�x1?�gG�j�\�x;X���\��gND�0*��w�6|Ŝ��aTњ�c���ЧJz^�~A�t��B�b��s���0�ɣ;8�kIs��*^�V�ObvyY����W�ߺ�0�;��)Q�/���y�N`j�m�p;�����v���u���i��DnX.�pKd��l{
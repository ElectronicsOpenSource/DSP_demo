XlxV65EB    67bd    1680�e��b����u�bոlS��Ӥ5?9*u�a=���
��4~}	~�T���ys�}���.�Qy��"�l�:9�x�ڭN�N�zf�z_ء��t���`{?�I�gZEp�o��qзe�^Y=ۚ�+I�u��6��T�C�j���S^Ǩ_
���_FZo ،R��k�80�g��<M��i���&��nm�Hd��v�>N�OL�g�ł��߄���	��mr+y�#��K���ӊ�F�&��7.>*1�
y��E�o��tD�R�A�3��"��_�/�t�CY���Pl[ۊ����˔�ck�8�[p�{�&�m6&�4P|aݨw؝v1e����;P�� ��͡���2&����$n$���|���'bΠ�W��(�(>���w+�����*����*I�&G�"!��&�/S�(�L+�.�^D��4��C�R���D�����&���������ݡJs��z5C�<Y�ʝg�E�(-)��lR��D�gS���c.��^�xks�$�ZO<� SxS������!�]_�Q�p��{i+<щ���,+L�A�����`���mMg����hí��
��tG2h���^X��|�I�xJ�
(ܲY���+�~o}=e&��U��rS����O��a\����/�EČ��e�f�K�\���s�z�q��ὼ�(���"���]��n�i�9/AG*�]�Zry����9R�Y\(U`�"u��{�W�8n]�=Hs��#5���@�M�O�Nj?�I/gN|��P��3n5��.f�GҖt�p2�i<��+����[!���]%��L�L.���~E��#��Q:�2RT4�߅����/Q����O�c�V�D@�L+��Վ��s��Bv+hx=0�{�gv#x7�G©|��U.�T�C�]\S�w��=�?DI�Zd�	�67b2Ck�2<������4�jjZ�q��)Wf�G����{wX��wu�row���j�Tj(��M�h�(�&o�!ţ������1��`��|���g�n��o��A��	BY��3�����6�OF��ͷx����`��M��x�LP��(������%=^�_DY��Lq�eJ\�Ə o �:��_��#\��1����|�r�ꢫ/�s,�XV��Ӳ�3<e^eBʶM$�`��:7���
L�5�dNѓ��������w��d��a?R׾���5voO���<�Y�)���c1����C ��ĂူF�/��}���[�De�p��oԊ������~���[*Dyř)�D�M�|�86��wуct햕������He¶����2��h2�mA7�c��=���t��Fpma�����l�*Ԋ�C ?yg�h,�B�[\9i�|��c:��r�����}an��AĜ���G�>�Ưg��4����Y�dR+ݘ��(3v�`�ނD�K.	O�'�E����y��D~������J�X��s�IH���)p��q5*���)���-s���6
M� �i���1cAeI�@U空�-2��<,�x�7�ڟ�<G��]ґ&��	\���� ����h�L���#��=���}E)�`5�f� iQ��R�%ȲI�'��</�<7��C@D���K�r�"/�Ka��-��o���`e�Z�"��N� '�x��Q�뇦� �7�o�K8(�򍩛o�$�gy�*%g�\x��*�ե<���Vb�H�~�24�{:���W�oK�N��Y'�&`0 ���k�7��TG�v��(M���� ��m�!��-X|62�#]o)�:k��X� φpp�����#!۩�(H������3dG�@�H�`O���0�
�6~��#���X��ڡR�����yWmM���_����G� &�f�
G����'D��ah�*
��$��|>��:��w��M�1�����*����F�M*���Ē�N#�x�<����N�����dLL$`�!���[��oH�#qH](���o��0W�-N��g�>��R��>`�������8��
ٍ��2���|3�X��
�{u˨�Җ�ti� �t��ିD����u���L)L2��ޑ��\��%N�!��il;� �lA�积,�C����h�V�v�_������-��@�����
�_��kn3D���]�aI6m������?� ���/��U�U��N��Ҷ��L c�u�>Oa-ڇ@�L�n?�!r�)���ϘM��u���(vS�]�,�Z�Շ�[Ain��R���:+R ���;��@0�!�c��4W9���o�F>�6lT�"�(���+s�ȡ�o�aA�J�Ê�+<�/���:��;ak}tŷ/�7�,�M���/�~uo��E����i=��Yp ��5>!���t*bӚ�0��7al ����҉Qk��u���Hn���N	*�{1�'L�ݤ9�
h�)�M���!H/��|=�jAF5���^CH*�Y�S���vڮ��C�#�����4פ�
^��%�f�$ GH�$֛���byZH�R�3E0m���~����G���Cc�*	�d|Q���{�a|�DP�>���Z��|3�������V8/w�o/�h�Z�E��(�5<T���>�N�j�a� ��{r=��S�o��@8�m�|o>>0������g?`�T���l����+��󩈑v�#��5L[��^��f	��\i��3�4&]���b0%���#U��/+R7�Y|�HN}!��Đ�����v�\b�Z
�O
8��}���T�i1L�gzgBQZ�\��E:ƙ��q�z�;��zY|�g��_�k�������tT��s&���}z��@����Co���I"�Rl�y�1Ew����p��ݻ_l=��@��G.�+=k}#��q�s����>BF�~����N�Hwm����͓ycu�m��Պ�25�o��B�aH3�ʶ��
�_�0��������p��Œ�V��0��d'�&w�������R��Di���(�R]e�R(�V�
s�#m�J&�`O���
<��&fxix�udV}״�z)k���iR̏CPi/�|rѿ��Y~?Ry�6J�KFĽ��z�H�$�v��	]�ᖗR�:�*���NDo��G�?���T��B�>	��ު�H��c	8�3@7s�|��kp�Z
]C@j��])]�uG[�?��#��#RGӣ5U�?�1���V�s�ﴟBl�<`٤6��o�l�,h�'J{��X��Yy=��zH@�Ď|�u[i���2��O�adՑ���;��.����}ϛ�D���P2�{8yA�L�>4��B�.�7�S�*�5V��T��$^מ\daj�6�M�#yY�X���KO��bۡ�;u,A�^�qL�8��ծC�ES�r��w�րX�����Y݇s�b_�=臽�.�ds�1a"+������ɪ�I������X�!�Qp�L�[�f?3W�dw��%�~��Q�@�����(�7%���z
%$&%��:DY<��4��u��{�6[��rJ0�y�1c�[h=���'`.&t:S��@�Um��zKQ�"�-rR�Ӏ�ls3h[�����bEiE���[�<�	F�����=v�	���#��~b�$�2F=�Ο�>�L��u�NQR3�\=��)N	a���1�4p6��u�S5�r�ι����m�<�l�תH��W/��pq}��y�y&k}8T7G)NnGF�����-�t��. ż#�č�H�R�����R�l<ˍ��<����G�&�����	}��[U�v�	��+�V�CY����@��{�7Z���Z��	�I"�c"o�8� X����V��)���hp�`��ޢ?���Q�$Lt|���=ީ�c��DTp!����X�љR��;n����L�'�yY�p}>>���b�x{���e+)y��9��şG=��6��tFc�E�ep
Q�>��KD�Z�(�Ĵ�
&���}����ڴp{�#@_���]r���_�w��X�k��j�{X�b�� mt������=��~�e�
Ba�L%���s	+�D�ݷDXױ��i��9G����-��Yi�w�N�{����8#Av����T�ݵ��;��(tυ��J�����Pȑ�ͧ|��^�1����"j��@��;�ka�sE��S�1��h���XWhp�b3z������@�J�8\"hȯ��@hp��iz�! `SRe�+������n����G��d�SU;�GQ�6:5s�ۙS�I�8��a6,*'mphGd ��cK�?��(�T���	���){
�"+�zd�h"���=��K��n-, �V�ևyCʘ�[7ks�釢`�Z�	��嵌�1͒���ѴT6����&ՠ��WW
cQ^=s���\ ��%X�LLƭ�x?�-��go�+���H�����3����_�AR����# ��}���3����Hrl�)-�[,o>��+���тě6�=ba�p��}Ы�D�1��h$X�ĸ�[���ŦG~��US`rt��sf�M�F�*B����c�d8?J'"#=(<%�gp�Y��V �gA,Rף�m���E�[�=�է�#,¼"�q����v"�Q� %'�;B=0e e�%C�d���,c�0�òј3"��>�'c]���3Z�����i�m�>�{[���m8	5sB�	�| 
 �Bd���cE��\��fA���P�E��8`9���ioz*v.��,X&!}�u#GF�MJ� =uZ�w�mh�P����"�e*��8$�x�O�cn̘�ob���c�I�K�7�� TN��@k �w�?��ԋ����XJ�(���	v��J��4�� ����� -�j<�P��4�B������Foꉯ�Ac���"���n�pڶ���Չq�G8T��^u�Xpv��(;���JA�3e N�J�j��47K�=����p|xf�S��4�UF~����] l�v|(g~s%U!�?�#j�� ��c����0.�{tD3<�0�Ywv�y����WH*�pf�'*���j��Y�����p6��)�<��FP��̟a.�<����ׇ��6p����kT� ���F����9]s1� �8H�L 39%Gz�^���ּ@�,4z��1�>�MD$�!�����**}N?�#�ICýFm8�D���[o,;��Z`GI4�Q 
��,0(t�+R`ˌ����|�;J+�*��bs���:������)��K���r�>����ZG�����g���'�w��,e�E�������K�|ŤR&e6������q#���
�t�T��i%3C������՚"<A��Չ2P� �x\�敨K� �\���Q�5*9M��x\P���.��K.y6E^tC� ��A6S�db"C���_jj�7)�7�8f6������m��Ҙ"�Ty���*=�Y���wyY ;V�{�x� ?����������q���O:'����zy,A����/FtCF��+Pc��"���+�cpu�q�����ݜ��\X{.\�p.���t\	j��t�*$b!�Z;�ǝ�gA~D6���	+8StA��c�9�;>���fp.��6�n�=���VU�|I��f�O�yޡ��d�{�=����/�
XlxV65EB    fa00    2fb0N���֥��L�p���U��9�C)�cF�QCs��<Y��	��z��w��1���Ð��}�R�1F��w�X˓����":1���{��X[E<ڻT� �Tş�&4��ܪ1��R��F��{��lc�d�S�Z-B9M|�w�o��L�^<����+�A�V����孏(��l֐�Jx�I mU��������^N�	���q���g��Y�3�!�E�קR~Bq	����HB���g?W�s1����O������`ǿ�r_��2��������n��S�ѧ�d(��.Mz|�3��"a����>$���ˁհl�O<ኚ|6�W��,�oK�2���+���x�o��=�o
����%�R�1�\N1Trh�	����m�.���PB�APȰ2���������t&�MD�{��;��C-�e ^�k�~aѕ�q>OuҤ�e}�Fk&�m�-��geb��^%�ΩUJ�8K;2+�շ���[���Q�n+�#�fC �B�&��`����Pp�tG�DEK��C˺n�u�FI�Ν%������	iO����\I��,����U��1:Su�/�?�
FȘ��.��@���l��N�?]"*Ҫ�H¹3�(��g��_�������]��*�x�h׶bm�M��/�h��y$��I��9�xP����Ǔ:��i���H���ڄ�W͢�&���EQɞtY�q��sA@xy�R9����x������=�Qy6��~}��#M
��FG����Y+�q#^JF�t���4�"TF�-��h7s���0:� L�޾���{�CG��zw/|��ow�D�10o�B �d���Z���fl���������$����Tc�Bֺ��SDr���&ޓ����~�O?���u����N@��~h��K��@�ѳ�n	��L�;q�}[K��e�	v���7f��T:pcҢ9H���am�$�LΗ��[�7����9��1��aVY��Ѳl����)������!�$���Ε�=�X7����d)+����9K ~�Ly/���'���ʪz�y�5�H%P��S5�,�.����l��͒ڬ�p��5nuV��X=0mUw%��Ӿ��ͥ�N���{0;5@9���x*	A��؝{0�K�t��gnV�W�
��Z����<Q<��;�!���>ù~W�J�z�C*�mi0�U���wP���.�MT��9�i�	<��Z, ����HǦ�������ON����� �ZfD���Ð�K�{�����|�V�����bK��,v1���o�ם�1)�����+M��\p�p�g��
"F{?�Q��)�Ja�L�(0�29�ۭ��T�_���{#?�N,CA'�^�b�=,.7*;?�c���^n�5�V3�Џw�>O�q�&���l�ٓB������X�	K�,J�=�LP�.������ӏk�mhX4U.-~����g�&��L��yTC��ͷ�P)�ܲ�h��"xcvAfG�gJ�-Ξ<"�"��uB�8��1���nGlY1�'@�!+��O�p�Pq���"�xR�����J����CE-2)$ʭJP=y�����ƻ'M�n3?(��錡j���k�JNԋ'�@��P��CG}�S�@�[@��_à��3��|�Ă5ਨ��z�]��T�z���+�*��4y������>�)y�����4)�:w�[��E�p���뼴1n�B�:�O�p��v�e�~[/3�-��_����y�?�@��cZ�Z8�h���^?���(�Z$W�z���Gwu���vet];���.
@7�Ǩ�]�<@ZA��_N��nI��.���S���h�G�!}�@�/�kB�X�=�d��{��]֗��O��#7=s��Rx��sb�|�G8WKa{9�dV�=ٹ�c�T�q�Lg_ 
�W�����2
�]ԑ�V3xn�.j~Y����M6�&q�$A�C�"�$�/����|�dQ/"\+q��1z<bu�NtAmuEN0�C,V@�T��.�c����<�0�Q��M�g�Hy�R�b�D]=? 
��$�� �������}��ݻ˘JW]U�N��z �ܭO�	��Sq����;����E��k:Ư��CK+ڈl4{���`�|�è���uh����XG�˷ {�#ب!��*ݭ�+KByv��-pi�\��U��ž{��<����)����~�+#*N��{Ŗ�1dW��HM}^6�>�������E�/+�����N�8��;�a9-�K��x����~l�[�^�pp��{^�W�e�c�༃��D����<�N�)�b���Ѣ,~v2G>�u�QG��0��Ā�rBx�0�M`���%ެ��i����σ�'  ��A7bW��
����|���Bi!:(�U����\��Ou������ �3´0S�p��+!�Q}Ҧ�5Ƶd���T0�>V���S72�2"j*�D��2�L��%Z�O���T��5�>L��o^
��^�n��\-G�!�O sW�LO��a��g��!G�� �k�%x4�}���4[h!n*G�hC�^]B~:.	~v쵤�$g`���Rh�^�_�\ū�0s�U��/(	�f��&Ҳ�b�xT�z�
j���QD��f�|c�׾$B��u�|�	ľ��m|��C[8��ڪd�^h���wY��t!�۷������#!�\q�8���_񯠚�$~��.�"YwΐE-S��%���h"o��$J�;Y�˴�i淶QB�� z��,�g9�i�᥃��"%%��A���L�w�NM��Ű���)	�'���n�_&Q�;�����ҟ9[|��k�����5�i�[������ �f/�]�������(S�:�3`�&ɢ��T��Ιq�5l�_w�S
��ԨkW{xhNG4������A>�SK|�d�?1d��T�����V[�H|�6M�v`گ}bY�~��U$LY�޲eGWg� Ҙ{�ZD�p��OM6u�9�u��L��0�]���@d���ӡ̴��%�0l��?�s�O`ю���>0���a����H{�-8d��	��1�EJ S�gK�`�!�e�ݕlP�`v�&�C�Tr� ���c�&)���p��#��י .���u��YG_�/^Qc���k��p�j�C����r:���"Yo#�zg�#�)`�)rk�u1tK���a�@�19=6�8#hA���8��oZ��i�&A̐ ��'�m�֮@C7��5-���|���
J+��[+�b`�,���&�+��3�J�`L��a�G��~��:x�$�_!�k�:�qf�5��E��m�4��Z����5�ӣo�@H�d�̃�S^t#9�P�Q\x��./�5��?��K��4`!̘����8`�Zx�#f�B��q�'1H�@�&�bbQ��^_d�+��wjE���[�9&h���u_�$"E����ic�"F����Ѣ
�wp�2Tح�Ϧ���r����j��\�h��N�r�0�]9ۮ7w�d���߭��*�s�i.�u����2
�b85����,��i%����o�]J��H%b���x�3\{5����Հ|�G��lm�_��e��)$�r�At�)L3��	�'\$E�[�w��r������3Ԙեʼ�Oޓ�L5D��F�	�q&ۿH,	[ �_(��y�S�C�Z�� ?�N����%Y�-ML9cn�	�I�^���q�P�c��ܴN�p�>bx�bN4 �.I�����N�Č���	cX�PW3�	�����?��غ3p��,��Hx4�U9�ӑ��s��վ��)Bn��Vt��v���g>K���Y cy97�f�ڛ��`è�Z;n��,���5�\��S���=E�u�Ɯr��JH
�A�h��\���ń�F��W��u�D-�a�����I!kF���=���sN7�xs���������,�b��#��P�»�����ȴ���D���|�z��Gҫ�&玑������vaq�+ ��/hAa0d��:uW�!�|��ZS�U���R/Z
:K�\C�+���J�RDU�{�g�����A�e�RB�(T¨a�x|;��mb�h�*|^v�/�e��KJ!Q\3��r�ò��L�em�Ȗ�Y����r�w�b
��A�r�m_�ȳ��ӯ�0���� ��	Ӵ+-yҡ�?�kD���D%���"�O�j��)�f�S�c�9\�(��S33)�b��F��x"~����e�z~��Q��\�Os�w�w;����+�����"U�H[�qs�ӵ�k��E��"`�W����_C��rr�,qclR���#~ܞ y�~n*I��\̽�}�i%W����2h4�e�U�s��J�a5������M�qڮ3�6�����}��;�G�Q(B���u�٣3��e�#E�~3�~�)��#�p��4�ŋ�#�%o�v������2��WV���Sna�̧T���7��m���;��ROK�! *u����'d�.N�ImN3�g�؀Fr䳿֌��d�%�SF����y$�PҨ�_h�fgYBCyw�My����N-��a�����v� ���V�mO��FO�<S�i.�� }�<�Aa���B�Gq;��|um�qY8�S�	��V~�P�Y6*����2��&Ɉ�:ז��)RI�>/Z��Ov�!O
r��Q���0VvF�c�h4�4R����n{�������]�5Sg��s0������l������s�� ���z�;��-ȹy�PB�����*�:aO$�G@�(	�JS�y��{�-��0�N�&��&jC����d�����c?,�O!�����7;����}-�|���n��.�!$#1fK����:m��iK�1IX(KO�������
A����&��s��x{noH�&C+(kX��0���kt����ܹ�U�S�X��pP�i,�ˀ_�m�ckk}_��F[���#�
�Q��_ �Y���4�
%|���%o� Q��G�lsB������#x�	ies�%�1�x�� R���G˘�0��]P��«Jh'a\��1��u�L�TW�\\�ԔFEߺ��<	b��� j�Ҧ��j�Შ�)���5�k]����R�=;u���)�<DM���nB���k$Mi7��������M$0��QC˪�\,�+뎚�H�E5��촾����Y[ǛBn�W�����-��l/�x�oX0|�.rӊ�dì9\3�����u}�[��H��S�4� p��\S�8�.?L5x.�J�y`1���i ������K2x� BH���qʖ}���rؔԬo���$����_�Y�aҾ�a���V!n8P�D���f�`cG�:�����HyI��d�	�I!ɶ��g��ٯ̚[� y�K�y��K�����V�������뮑eu)�;GpAR���A l���	�:G��:�t��51q}�~K�q�2B�@Tjn��3����հ����������=d�~�Bj���j�3�Ƕ-b!�8Г���u��BwD�5�����5��D����BS�$��n���p��ߢ�P��t�t0.�t�rq�S��R�?��nxS᭬ΆUVo �M�MV�1�����įY%y%?<��7V�B57K�(+�X�rz���,����s1���.���!W^���j�/�-`��=X���}��_��
%7�߱)o�h�M��7��?�͆�]�>�3Z&����ν+�D7s<��>�����5,U�cg��O;iء�$�_����.Z�4RIᐮ�h;?dw��`�`���������������Wj���rD: FX]>�s@��3�D{�St�=93e���Yr��e��&��#���M:����/l"�����8��& _3
�G�xȕ;�W�����;yw�̍�T�RP����kl��\7|p:�-��b�������xQ©D��	���8�h��h�-ߣ�C�,�]��W#W�m�8���Ǌ�/{������l��]����d�$#F1�q�1'P։*���Ә�k�Mz+��8��I�G\��z���GѾ�^����=�{�o�e~6���U�-���(�U�;W+�1�ߨz��'E;���Ӈ zZF����4�{$�C�̚dM�9�e�ɩN����7e[�5ʎ�ѹݤ���{=��vƘ��mQY	��"a��so�z犅\�yj�2��@�[�SW�^|�d�jŽ������M��U�eP2�N�^�0���\mĀ���RG�A�5��K9�9f�&�!����$���e�' ���2W�j���46q���Zn�|���EP�Թ  ^��+ut4hq�����|N�W��0��f�QW��rt8�9๯ ��S0��v�kps��w����g8_W<9o'MΡ���+ǗQp��~,�w���H�,R�$�8,Wԛ.�ɻ�X
�L'O�Tw����JQ�&ֶz�pkZ=���K��䲇tth���z�
�m��]���#�t�[c*�Bb�n��o�)s���ۍL�	5>g�4���� �d�k��;$��[I��v���Vv:�7 3���%
"�㚤�FL�pIn.4���p�Rwi	v���v���Td�*r����<!��`��g�.C�+HH)�^�Y4BZ���+�`�J��ތŔ�2%)}u����d-�
��,m&���6��������p_!���(�o��U�nn���D*Z�����kvw��â��
�j�IB�P��dv{&��=����`V�#R;m���yAcj �g �����ɼ!��O�t�Ƈ}�n�I�:��!��?��	�>Q�	%�s�	ޏ��ߞ/�����Z��Jp��W�'i.R�����>��~�abv���g�X���(�I�������D�}ܟ�'�&'�X�_�5��mEC*���0���Y ��g6U���C��C֭�'2]&�
�;6����#o?����և!ԡ^�;X����	�����u���"m�N�;�|5[6D�N5�̐�lJ-@�e��n�K�k�(�+Zș���ox���jF3 ��˪��d���}��{]-�hH/H2�����a;��w�k|,D�3��Wz)��%��JO�����a���Z��IawB� ��X5nxL��6,}rD�Ulv��C�ݬ���CE4u�,P}�-�& ��1/#�Qr���o�d����t�t�3���љ��]���\9�G�3_'��K)Ơ�op���ʅ0
�&4yP
\�%R�b	��y��(V�0��r�r�d�_�W����dH)<��x16�1�v�K���v6��r�̈́k౅-焖&=ݕ:?���̒,Z���3V/�Lp�̄�.Z"���#<�1E�,Cİ��pR�"8�-���4`�I���ؓo�*�4��ه3ә"��W�����8Y�������f�Q�z#�v�[��~��`�z�1����JV<���$.Y�)��Ǘ��$#��'Bf ]27�~-C>uX(��HgiQF��e��u�H�إ*G�I�Ĕ��:y5��"�W*9D*9��.}����GD-M�?�3�/�AC��7�i�F��� �~4	А�Ye<.�t�f4`K�H�����L��'��\������6.@�K�����]^���,mr��8ԡf��X����������4�KJl��Cq�\uQQk�M�0uh�J�
Y���:�9���,���Ծ̏o��A#�����bϫ�S/bw��$X��C��k%@�nB�W��ɛ���b��X�}?�	d
���>���Re)����n.Q�B�1�n[�?�K�tZ:X+|�ߤ@�G��I%0��E1�h�����/[�Kn����fN�J6PE�<mH ���Ŷk��R1�T�(�T)
�S&�2�;�s���f�e���>=�u�����lRC{V5�N@��<�^/�eO�C_����u9%�h{������I!�a{J�][����<F?�[z��z3���O
�ϋ�'�e�;UI��1u��T��K`�f�����iĺM�bY�9ߓy���(��I�P�g�)�����Sc��
Bq��כ��R�B�����ٙ���+�4g������'��u���6��ǟ����$=��^����}��g�#�EN�e�\�DD~m�aN�gݱ�e|"��w�z����	˷�T��g��	�n��?��^.n���]�7�܊TO�sǆα.�,j���B�7��-mC�#n���ƒ�f��Y�SdNu�w�`��ز:9X�-�i6[�`�t�y���q!{$X����+�c.cӉJ�>����͵���	/�p�O�w����r�S}���0�)P�X2�"p�
�w��i\��ߩe����L�PL
2�.ES������U���B#�L�Q6�2�y�+,�ߣ���,���F)DL�d!J�T�׎K���!|��VU���\H9G.ʔ�=j\� l��x���@�o���%x$�=�B
����s �Ac��� ��P��CL����$��	�I� �K�����h�囹���`.U�n�f�������Hq���� ##[n�⥷ ��q�.w�u�+�_�Eg4\�n!6ɉ��a�D��LE�</f�7�}N4�OϽ��̓�͘�,��z{bR���T���o����x\���^��o(�~�mF�>����%�M}�Ef�}^��%�O.v�!k�G�Ks<��_i7�"Q���t�a��(��"8�����_��5 �ZZ���@$����D��=�0�H��G�P�����g�;�IZ���ϱz�GK�U�h�+����26���>�zх�RP`�$���,�9Uk쭝�CmB��ѪՆ�0���k�����`M��İ�F���O�gn��.��^D�<������u��<PB��n2s˘�g��L��hNq�˳1�mf��N$�y
�����P��MG���E&'R&�,�d��^��H�}�l#M��X�'+Ћ��):w���ןy���n� i�1��U.Uvܼ�\I���8�]���|���r�Sa>�<o����o�f�b�t5E����w���Rҏ�5�>T�%��A�� �K���y����*2� 74��%�5�a�~�,t�9u���"����!�w����!7[@O�6������+E;E$)i��M���М�u�܇���c���?��A�iY����k9�@d��`'�[�Ce&�q��qT�%VG0��=�,٬]=n����W��-=ig9�):>"�s�$.����gNu�L*x���z�5�j}�A�a��Õ�w���"u�xϸ��
=�/�_�t�k�J=B<E�-�(�m�}TS"u�J*��X P���7���]��z�a,z���k`'�]�ҙJ��3��ݠڀ$7�㰨Fn6�4���n��+�v.�s߁�D	��~	�9`~�	�ŏ���\�� ��&߸S��Mz�j�p=�6Wsk��V�_�|
�ܖb}���A��)�
>?O�ך����h�G J���)C}���jKj8:��z"��\5^��&bd��%��8� XCY]Z6�ѪE��:;�`B���)H�����8j����'Y�,��������(����Q���n������,L��p<��N�� [�S�}����H;5Vw�ӆ�M7A}�\z�D��i���z��2�.��DqTk�I�h�����wa{#B���X�Ҽ����Z�B����M���qP�t2�h�ޒ/�ĆIU��@Dbʄ�hxXW?����ς���٬+�l�#D�g��|��4t��%�naJ��ᖏ����L���޴���<��Ys��
n�����4<�; ���e'_��*�B#�i������و��K͵��P��~��{w	���7��%(d����
ppn���F�����d��VK�Q�@Wv'B�1�x[��>ǥ����f���Tu�Ψ1��5���A�%&`��8��;@�) �xM:���g���Pi�ez=�0��1`x�s�����·�_��[ ���|�VR��ez D���M ��exc+�,]bsC��3>H.6V'= �W@���>�����!�]nSO�'����h�8G�{6��p��N �s��ܭ/��*0S[o��ff�,�v�/���F�~�Ɗ˓�a2��'� �c�*��8G ���*m� &�R��ں����	:>7�#(N�"4��gmG:�{�\����X[P�����l���qt��Y���I@_�:������Ò��b�K����׶*��qL�[b��ЂPx�|"�L�y�-��52����Wݠw4�2\h�l��d+l��_����ɽ3"��gBn-X�o��X���~�R��
��^���S#�;��Ɗ�k�"�ޔP.
��A����v�\�O�UZ�:�4��ա�w���0F�_3��q�e�7��>�	�
x6J/Y��H��e��*?�h�,WX\]�l�F#��w!d����j�����kș<�^��+�G��{O/��	��%�U�`���#�C��J������T�|_���L����Er��j�؁�\�Oi��ue�4��Gw�i�	Y-���c�������ļ�ڱ�*F�6� 5V�l�c��Ox��n�Uj���q��ֈ�qp�����6�`��g���eR`&�!� W������gE�{�[�9r��B&=�Ǧ�;��P�� ��6�7֬��F!9�֚������A��S%X�!^�:1���;���r(�N�/?�)�����4�~ge���q�h
ƨ�y�br3�t��z���R��c]����
QU�%�����ų��h��������p���c.�A�t��n6������Mǐ����I�"��+L9�V�n��C��OOr�u�7-�FAǉТH�c���Jʌ���t��E�fw��!��@�v`d�H��N7&e�	��GY4�$�c�)�>�����Vo�|��\2��s�x��R펭a�P���-���Y�\���\Tr�H n��c���|Pr��cQj
�����{���կnW�Ƥt�;E���1��J12ӆ�B.x^�����yX�\��U5�)���5�`���xI��
� 9�"Pه�2C�5t�|L83D�4�[��f��Kp�y���_����Q}������X�B/��/�0�����i[=�j���=�N���O[���D�J��1�6�S��)���.�KІ���S����)��;*�19�#�3d%����?E5�!�V�u�������Vh�)�r��^df�h���"�����p�/q��u�� �����)�.B�4�O��K4>�T��S�Fʠ},�F��>k�<
[e�0�����#v֠����3c�&1��sޯ2�.Z�0t]��3V=θ��&1�����I�_yr/��"~)nR�7�j�[fw�U�9͎�� ��d���RR\"gGd�/����'�+�,�S�=���F����|�3��O��)ZE�-����F���.��|��|kc�չp)��}�����#�o��׋6>W���X<� �Th}��]�R��NE٣Ȥyju~I~�gOL���ݘ�5^��4a?�؃��L�:L�/s�eR9��7��ƴ~��h��#
�����pYˉXⴓ�]�7�9��8zAk)�jxטA�4Í�!v�zw�_��
Z��9g�7���O�Nsܒ{-�U�cA�RqoA�*����i�Ǿ��̞��Lt�%+��q�T��*-�/Ji-��k\�t={!������!���ct=I�9̕m䟃�B �]���;��H����x�5S+��)&��r�%�C�o�u�OՅ@��C��;	�"ę;ZA������Y���v`�l�s{���!���JR�BCcF�2��7��V\dYꃷvn��Sq�  yp�nA�Q;ʼ����ߥ����S�aG�f���W�Lҩa$�mԄ�V��CI:���.�}�{��0�b�j�A�"�C<�]��?�A��Ą��DRO4d�t�?0���%�Op݊ؗ�V�l0��7�%;3FyQd�����4ۦ�HyG��g��
tO�ƽ=��֨��w�XlxV65EB    bfbd    21b0�gҍR�*���|~2O�%]�eǍ������ސ��c D~�A��0�n�_Π��}S>ʫ)��0����M�_��� ʵ�U�q�M��|+����#���Nd(�1���.��C`r��k�-�l��$^��H�D��ԔL�.��_����s�|g���*���ܷ��s����*�3,�:�,�P���l�n�/�o��ɸQqn�\T�- W�l���Y����<���IlZ�������+�W�dG�RfU��ͤ�gk�Gʔ��Y ����ԭ�������1ѕi���b���pn;oZA�u	�g��d��FHo ������"��{u6~�H����э~EWśc����yw�G�f࿊���r���Q�V�+ жDЛB���G!$FL�E
��?��nYfW͵�ֽ��#�nt�V�]���A<I!M�s���܇���ʾyr�,��Pb���&����!Z��ׯ�bK��-�i� �3�@o��喾o[��ϙX�t�(���YF�;�|��@���Eeu<�ɔ9�#n@��7QN��U@���j�7�y�pk��MW%����7G-���רˋ�b��X6�sO@��Z��JbF�
��B�	49�dNˏ�0�_;����e�������=�4�q��_(C�7��P@.a���2\����(���P��JoE<�R���l�$�_я
��A낪]6�#I�� �B�5�üg��]C�}V�Ҕ�#V��9+C�z�Q��j���c��r!j�Q�<пm$2�O%3gn��6k���/�Q�_?�p��#{^�y���ٖ�T�m�jy[ J�i�hۮm���e2��z�)��a4pd��7\L�q>�f1�e�K�/[����k�`7j���������i��xl0��*H9 �B�̔g=��)O��ۥ�P��%>�[�%�ß��X�ϙ��B�	'U�Fm�\�?֗>�N���^������(�������Q�94�G�	q�'a��Z%n����N'�&ȉR}��@'{�𪍲��^4S���Ё:r�fG<��i�Ɗ����:~��vC���} ���;��01���Oi����3�&ҵE��YC[�����n����r>6^�p{8��p�9�v��lf��J�rHƎ��qnk,O�i�{���Q
���������݊�i���=ta΄*�(������ֵ~y!Ƌ�X�ȁ!
<���{M;����Z�l�V���!?��d�d���K����_������P�sC�����Wj���=T(�`��,G�m5��I�m+T2��,q��X.�l�Ch�;D�
�p:�1u{����T(�P�0��F�@���?ko�;rT.jt�Z���ڮC��Y�Cۑ����\�%�Y��	�s7�F��ޛ|��ĦRZ�)<\E杓S�6O̕c	�K:оo8���|����{���F�j�2��H����	��
Rr%�?�X����S���7a�G�(W}УdT�x�e�V�r�1ek��5s/cT�S	�Y��2ó�c1%Hz�� ޕ�%��F{Zp�ɓ�C� ��1�ʽ�>gY;�6�+%�&��n= ��t�&j�j�y���Oo���3w(+@f�;��IԤ��q�Sx�oF� $������l�-<!U�9~�q��i�ދ��<Q�Y��H����f!�\���X]���-�c�ez��|�%�F��̝�(c�����n�k�۶H��*���ŵ�(ց���_��|�eh ��׭�<����2M��aA���|2B�C�����`�R���E�����ZJϬ���$�(��/�l��~#T�m�b�_� U�ʅ~��
e����]�L�7V�%"j�)*�P��cM3n�$@�9�!L���������!�Q,�vsZo����W��C``��kE� ~��u���K��k�D;!
�t����e��BtQ!%���^��!i|I�De�v�/г��D�V�_����.�إ�.��k��J���A�l���4z����֌}��g�B��|	M���z��D�g�Z[����e�i=W��N�P��a#"62���2�h7�OKͧ�����I�S� �Xм�u=�͉\��vG��� M��6�� ��W�uf��E�m�`��ۨҡsSs�׷�KY�x�qk��N�ؒ���u;�E0�R�CNbU�"�#鵳ou��;eg��	�����_��H�o(��H�ԍ$��0˦e�B��`��= ������%sƒv��"c�߮�3D��?��x��'�W%�H�Q���}�3��dshy�|��
��$���N+����0vӘ¯<���}��׀��]q�w����qܺc�~'��0�A�ƾ��  -�=���w�N���M3reF���<E(��v���]��e���9��e�������C���[y��k�:�-D���%�B�b��CX��ߋJUy��	�C���m�W�[J�N�!��^�5J��/��`�i�VjGh�֗�҄I8�8�"Q���˫�r�o��� ��E����HF��%�����U���[�G�"�
Pe��E�I9�*��^u�uok�=Sl�Z]����;yR��=C<���B&n���~y��X&�#�#���|q6�:yǄ:,#Rs�� ����c��w8\t��f�7�Y*����=֪bV�K���i;d�O��D�3�4!�����i�,Q����C�?��g����fd�r	���N�����fP�>�5�<���s9]���)�ݹi���NݿY��gW�Y�zB��ĸ��+�&�����f^�5(�l:�~=c<:�;|+�̯-^ʤ
�g��i���O�ùa������&c���ԃ�֧�#&��h�Q�*���x0.9��S�p�����Z˟o_�ԏWE��2��Ч�����|�+�������Ƅ�J}^�G٧"ߓ��`?���+~j���a'�*�hlh�	z8�����S�u�N�W"iu�F�g,��r#rT�k����@���X�b���Mj�����TÁ ��P4�7����ܿ �.̑�xdb7'q`e���{�o�佡}YA"� �Ե����k�:�DԈRh��eke �yN����D>8��+}uf�b�U�Z�!��-`�,�(D��1��C/a�q:��m�>�yZf3�ɲ�;
�O;9�-�ص-  ���$&O���U��僨�֗'�|?�MI�8h�{�(bԉ�����Ms2!&���+��'T5����H����3��!��6��PH��e�YJ��4o2-�@�b���T�t�|=4�ڜM�����nQ�
�_>�����5Dј�d�e�ӈ�cq�����<
���A|�у�/N�Z�X�V��^[�0���tJP��N8L������Ks���kQ~�=~⥡O��$+�a����TF��|��*�����������L���%7x����{0�zBS����H��&Flܻ�6��(�U%x����{B9�L�z��6�U)�M,�����=-&x�	~Gm�=�� �9U.�|([LCG���l =�J�k�c�!ONzt���H=hM�?Z)}�JQF��h�,�o19+�۱�u��_q��
I܆km�約����H�Y� `�F���i�(IHNu{�ѻ�0��S]`+r�j�a��J��zSx�������Y������ꃿ�%������M@[f�ydt�C�ȣ�d�[�bdU澱�I�4+�e<zp����(��i�g�B& ��6Dj�+�@Dp/�A����������˝�i�f�U4�Ȕ��aT��|�E��[p���lg�8�0�|�g��~csWI_��=�c��[����]n¾�:T��X��^)R_������KD�0h'��4�_iE�~�`Nsd���	��e��	�� ���$�B�q�2�|��x�<�pl(X�76^�l<*���4��C��Əj��:|S�CP���*�H� B���B��d���-V��`Ր�?����7_��%����r�z�����7c�WI�'/�;�_>����c+S��v&��X�wHO��R�D{�}<\� �_7��N��i]k�6�љ���@�����f$VZߝ����,�%�1 ��$Sn<�4j.�q�V
��U3�:�R�-Q��*�	�9uG���������99~�,�7srҼ�n����R�N_�ݐ�f��T^C�}�4��{\��k�FǄ@Ƨ�bòA.Υ[A�����\����\J�-�U��*�!l<��
�:���7�'�_1�v�*�f�*ʔܯ+�N��_��QDE���@a�����k0/�c��ޮɅ�-�X4���%�=��ҥ&K��,����6�S���e��)cK?r�O��9<�q�#�(`�i-�ͻ�?�OP�+�3�e[s�m�h? �����Gf��ae3���aI䈅�&ˠ��Y�~ɢ@�@��Q�U�B/�֝.+x�jYi�k����Kaa��37c E��r�+,�s/�����N|����纯�6z�Yǜ����6Q	���g왙�h
ܽX���F�K�ڛ�|9�{i���/=Xf��w��F��r���T��.q�M_�L0+��G4��#���I�`�4�5��(T�G�e�s.]���tu@a���3�]/�!`�p�)� k�ܼ�fWr ��{��7���>�Z}��=ND@�� �0NHC�)��%���F]x����������0 aJ�Ԟ�����[h���|im_0��*��s�
����Ռ3��Js�ļ}Vw�	����p�-�c\�zЂD�c5��e.{xۡ�����ǐ��Q���N=�q��
����8�����c��j�5"y)��(k@��*,��-�����e��8ݯ��7JD9��Z���"p�OTY��b�Hh�h�N��:�4�ձ�a0�/t[��+ըv��Z{��{f�G��
������~:���3��`J�߳�K�V2�,�ۏ3O.����!��֫}�zI�>A+�Ժ	O�PF��0�C#..��8򎐇>%�%�eK���rT�кC�1�K��b:/<��Ӽɿ���2=��'Zp&���`�p�ň���+h$Ĝi�
�gqD�NiO�C(O�����[�$�U:V5Rض�n|1>6�.�5�\H���9�gf�uF)%\MT���4os��\�cAW� ��Z
0�q��~y ����и�,b�pn��D��9rD���J�r�����CSl;c�t�8>��oG��o?[V�`��4��
�`"�DU�K��P@bƁ�SkR�Zl$!���ņ��a<d�<���K�NA�dT�M�N��ѪPW�,7��+�M��,�8�sF�Bh5�Q���~��������ev$m|�ش�Q� C*��c�D��GdC���2�a4{�}�Yʗ^P�޺�j���4�xgrn��{l+Z[C�E�|�#�8@�>r ��^���ƌe�)C�NC@冬�WL�v�1_��z���#�W���v*.��Q��.h02`���qJ5�>f�#�� �� r$�Co�7�eIȊ �(����g^Rp�	vv�j%�c� ��`�ה#j}��M��Ӑ��S)���9�Ȏ�h�D\U_�ǳ��zg���L^�5 ��-B/GG��듨�hs2B̡�n�o�XeCc5x/	��K7if�O�����_����'�_B����:��!ֈj�WX���'D=���ww ϟ�ez�Q��,,\���X�?���|�:�V��H���2����dg8��r�?���P�Mh��J��ZFU܂��f0�' �B��%�O.	�>�!���N�W}IA���ٿ	�}hY�-�6Ӻ��<�����%�H�.������X�@���ܼe�.��n�}����F�^8��&/�Z�Ā[�k]_��(�=���['�����c-�9��e���'M��\I�d�M��L����m6�6$J?�)~���$=8��Ef?�?a4�x������ �q#��4&��h��t����{\3��04{��� dڵqlA%�� ?iO���	R����D��)q�Re/�)$���T��=(�}H^H��_�Rߕ�^�	=�K/�uy;���c@'g!�]%cD��lG�#] w�`�d����y��p�T�K�gBF�H�ju��'���+T{Ja����-���&�4w�t(A�X��zH@�f���hn�g�D$X�R��ܯU����IV+�䦲��;\(�)��<3ZE'�&JKv��Oj]ۤ	)˚4?jָ�N���+qa�j��	��s���~�:�	O�����"�MXJ�SM6�~���F2o�ɠ����L�A�tGwKޠǑX���q��B-�$Q���� [x6�g�ho��ȴ����#��X	/����L��?�Z��<��Y2�]0�zVe��ʁ���q���w���#�&�[&P�_H4����Z��c�D\�ؔ����<��0ߍ��FC`a[ݤM�}]
�r�H�O���f~�>Ð���a��@�6��x�@-�cb��io+��&��B�n�U�=���`�hz�c�2�62Z�����*���6�O�8��⪡�e$Rj�Y�WTs���	��Z����,����kR��{[���K�k�p�˘fl�N��8Ci��Y��=$�&� ���l�V��٩�/�>X����b��
 �H�yg&2/O[zct�U%��W�
˳
mxŎm��|1RW��m��ޜ��{U����h�n��oF��m;iT͖�rm"Ժ=�t�lŲG$������ڥ�U�<E#X�ɧ�Jcs�k�"M��W���D���J�AcpC�u�Ӵ�j$�Vf�,JG@��?L�� i�릳G�J���[�n�ץ�0��]#q@�)1�0Nm�i_{U_����~���
����|Cב2�繷��9�(H됬t0�g�*�*��޴�G�9#fU�Izߕ3����F5<V�@"�,#������.4㷳$����;�X:emn��w���c�����	�H�wC��(���})	�@�^Pc�e�H��
��I3ϐ|*���^O'P�氥f7�����5��}~�~����B��8a���!�b�:y����H�é/����rei�p�6U��_8Ǣ�/�/�݆�����+N4�
G�.��'��b����;��K��䙨A��,5��
�H]CZu.h �[C��^�a�AC;ޫ��G);�\�v�Q������+%�lݘ-�a�S��V��zRQV���A�A(�m����Bs4-U�3�w�1�����:��\g������XZQ�i��!L�8kP �]
���)e�r;��W�b[0�՜Nt�,&WU$	��K92o
���n{��(�c^Z��კJ�Or��&�St\A��O��-!��&���)�0KFZ�ͯf"� G }�8mC�邶Wx�>�j�z\j�����'��)����!Bl�����~Ka��$�h#m�lex9c���Wu�qă�ݬc�w#��b�;�4��SD"嬼@,-�fI7�J~��o�H)0I��.�-!&c�(�r�8���Hme��������q�fš�=~��|��V��`�16h���
~��B(X'���攙��</71�}��:/�z>VO�w��+�}�O��7Y�6��>\.
9�%�a�hhr�./z<��`��G������*FI�22��Q)�'����*��H�;�h���<�CO+�r�ѝ�S��1$8`�QS�oB���r��:Z"0â*$:c�`���Cư;���¶�S4�|x��v��ޱ$��P4����B��~���9S�87B5/���=��zv3���Sk��e��dOG���^ ���ZO��:��_�S'� h~~?�W�t	6��� "}��y<�`��$a`�cl:B2^�'�-���0Q'D$L����#�<���px���&�����^����گ�[���.~�u��.h�v�L�����|}�'Z��YD<��p���Jo��7�m�97v���h�~��o(��}�^JVrO��g�����&�'�r@��Ȼ$?¢��ϭ�k�P������ b�'~�lA:x�Gu0�p���i����;��?By"=�r�7o�^Y�o�G�w�lӇ�I�$N %t���Oʕ1�'XA��6�F���v���}�F�/P#gBHR��g�I7{ph�p^���j@8�0zKdZ��a4�8E\���L#��A���0���S�g*>s����`�娱q����.00ռ�c*���T��ڀ�k	��^���AN?�\�ĩ�#��� �.�A��ùV�Q0�U����MN�[S�W��n�����]0Ю$V��埈��;@@Z�`Z���ۢ�ܠd�O%���稬�f<�a�����R���K���[���\+�qoV2-��1�B�������������͚�vFI�
�N�K)jjm,�䤲���
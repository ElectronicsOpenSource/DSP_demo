XlxV65EB    fa00    2ea02�)r�?|�z���a�𷃝�)�z�h�<�,+��x�|
U���1!�߉p�4)�IK�v7�{:�����^?�>6��sU��"Ϗj�Ĭ�LB�C�-��tI8+,�e�<)��aaC~�IЀk���5r���^�	q�.��=����!�*J-#G���V���%���L�'�p�(7�����2�梪��HqJ����T�L�]B%��%�y��+菌 iRUQ�Ԅ��ױ���#���{y��/���þ��vs�ݯ�ts��R����*��}���`�H��!��Ͷ�����}�LeF��mW|�*j豗D��t��BJ�:J��z����G|��v˴�[�su�4,�Y�!���d-��^p>�kb���iG�;rG�A��\�Ձ�T��	�K�̻�3��d^�Z"" �E��X�n祖��9�jGP�b$ʂ��}��rKhv-�b���:��O-����X�p�DЙ��[���a4�mؚ�n!w�z��TY~��6�uD�����S��v�6�,Sk�>SpU�?L�$u�K�ǜ&�l���^�}#�@K]OP�[�35!l%�<s��PG�p�xm��e��J#�3�oV�U��y�C�E����D^U���g��p{T"�J1�Pm5�AG�r��-hh�y�y��\�ؽ5�|���8}PM��	���������{N���E -]�� -ݶ���� O��iwy��W��	��M�,5�^����,�#%�ȒC�QE��e&�&�Q&����8VD�`T���3HB�[��5i�)ύ�u�޸2r�n�M�
2�~��(��grL�6ՏChk����dw`Nb��-�DشZ�׼�[��؛Pf\T��4��_l�W��9�8��f�4�e�o��X��g{�,�?�	�����l�ϭ�U}�Z�맔m��r��	]$��Y�f(7��+�����<�Yg�E?�������G���6$�ZC�G`Ū��}] ެ�_%Ma�)	��_�'5�qաDr�x0���
������ƕ5�1OQD�u����&�0�+cl����J:'g,P�.��0�\��	�Hi�2G3�ǁEM$]g�h3���e؈_R�o����@1	b��h���Oz�5�Si�z��*���hK��Lm��T����������=� ���r)�+�1�ܝ��Ls�#�ցF��\hj�/r���o�8	q?��n����+�s��4�X�m�J�`�k�S�Ѥ�S}��	P�1�A���Rɯ³zAe;`>KQ�b�Z�^�����7�
A|�c�%v-0g�]�u	�U�A�;nK��5�"���OV&X���0i@�B�F����4�o������*Ig`�j�<�����&�t��);1!��kq�m���;�b�/���	�϶��Oz�H���$`ۮqI�Jc�P�l��?��2���(Y�ǥz�$��4�c��\�ϝUg���=QTS9�᥎.x��C��=�*�炍�e7��t?���Bb�ցޢ�\H�o�ޑ*����H������KMG@��5<G�}c	[r+�g���,���0�;^cێ�"���8�q�(��tǶ��6*-���
�@h���.��p*��m6�K+�����Ah�z�\����{����խ��\�/bA�J2|/��M�� �k۴�o�r5#�Y/��S�M	����78��Đu*M���[��Ŵ	k�.��y]%��\���;�� ��<�oʺR�=��Hfp��k<���	�O���W{9����`�����N���QϤ7�T�N<:)Yq��W�]*_�j^�uUU��:�v@ᶛ�����4K#3)�@P�6�{Ǝ�l�����B���zu]˜���_RW\T�|����R:0���V`<�&��@�3[ T��{���P��7��+�tr��$�^��ZG�����^����i��?�R���t\� <��Y��K.]���?�)�����k*?���M8���,��	�m�x���jaA�A�����<��H�kƞ�l-�XɊ�a�%�
�����s�W �8P�`20��Z˸�
6oT�br�]<�C�v�E�ņ9�߲�]A���C�:������~�q�^�*��j�a�R�u�����IK;���|Uo������4ZC�a	ı���W|(�ޗM䢝� ����(V\������u�o�	��6�G�"	�Y(�@���a��h��ٿ�ʣF�hU��:��`ƽ�1��*i�HB��.��s�5A֊Eb�� c���3
�!������X2T����J?��Yh^�M�?F.�h>&��1�O1W�P��i����� z�Fŋ~y0P�B����8��N/YOXj$W��B��-j�TÓ�j5��-���*���*�a$k?�p����6�����eF�E���/�� S�7)�W�v~���p�������k,=}�Cdc�l琼����)ւ={8��a#�6hK�lk]�߁�y:7Xvg�*�;�1rN���Ϟ\���^�2cT��&����NieiTϼ�f7��kL�$���Ir"o0���5{.pyґ/�D��2�Y�����v�~W�WY��#Qe�?�Q��*�<�
�i���h������
!i�Fdd�G<r����w�o�@��-�.Bm:���e�Px�F-��.h_�sdbW�.�@��F+j��,��N5���5?b���� (����>��7M�Q�J������9�.��kn�l�g�
����H^ �_�C���S�"����^ſ�!AT�AA�C��_���[�D��$!�s����H�<�b��=��k4(��aH��ݭ��Y�m9��W��w*�5ʯ�>�kr�m������B����aG�\%��5<u:F���n�&�<:�򯎛�p��\�B��V�)��v�z�xo����,��kue4R23���^�\�f�CК�::�}|��ݱ���.?W��>���-H%�� �i�L��Ƣ�\}����HW��kU�L��p3�F�\<��TE��U,�C�����xZ�Կ.gը 4@�����GL�'3d�Bɼ�$��B*�F_@��쯉r<���ή���[h*G��ʣ��#ae4�G�1jK ��C��)��f�ct��8�晴x?Yо��ȃ�U�=��7b�"m�n1��:yŽm!ݫ���*X_M }�_�ٮ�H�g|����GQ�Y�z.�,E�" D��/����w�L���'4u�[,����W���K����z'U���瞄�.����E����i|�Uȸ�V�L��谏n8+�s���f]�T����~���x������P��, ^Alj��H���G�̏�=C0�aX�B�?UZϱu"�0֜c�mJh� ZW�I%dj"n��,,�
�=�,�n&��e�U�;i,���n?�"8Y�P� �������֞.Ϝ�� ��
�%5��P� zŞn�Ύ��R�Ԓ��жbWiR&>�osF>U�'k5�U�9���-B�q����;e�?O���lV����{�рɴ�E�E���h��Rr��>�hC#�dW�i���y��zg�@�
!��m*c�$$3��T
�6��e'+گ�H��&o�E���2��`t�`S0�v��T!��7{��c~>T�r�Pi�kF�X��
�����{_�����?��;RJ=�ww=��4ơ��~�|F�?�wE���V>Hod��3g��Hv|B��k�YY�)	bVsg��w�<�oI���c��ʼn�O�������
�wW`I����I3�f����#)q�d��-���� ��Ŵ�s��R�FM��Y�?�����g�`<炎t_��BV�n9�C�p��1���:7"s�{���;	�&	�'e�N�P��פ?�v��b�a,�����0�%D�&3�E7�-�a Z�ɺ��H] ����}]�q����,�Jt�H	i��������Q���ى@��n�pVzcG��W\ڟ�1�FY��$aAPu���q��I1 ����$�_bayXx<2���Qlx��;����[��rC�t1��,R<X�C��4}��mؖ:�s�,sQ�0��O�Ki_�Ʌe�Z�r�������RN5Ѵ���U7�'�±_��Z*Z-,�s�,s�6v,69zu"���W<6�g��M*���m ;p�+d�8��Rn��.��АE˭5��{"���L4B��_�/ش>6~�x�]iT�i�����5��Lt¯��[�6�_O�KP�n�����M��o�>m�s6���B���@�B&D.�$��J?�*����O,� f/p�%��H���^OZH��.DB�~��<v���R�?��"z�>�Iw;I׆�~2�2��P����dD4?b9!�0�Rq�����N�1VIxbQ�R����բ�;��VZ��q�q���?�^�R��l��i��EN3[�U\�ml�؈3���a#$��a=��dOG�r�ɉdTLJq��K�H�S����8�X�vٽ�oU�~]��GR�����ֲ��(*2���HGH�
_��!i"�i+��w�'�<��v�aYat�NO�O&�ׄ�.:%��|�� K�C�ږ��δ�m���m� �Z��~}܋�t��jim�ً�����F�Ʋ��)M���"2���FX͈lC��٢��nؽؕ�C����<���oWv*(N�����+�� ��dS�O�]N�2�����Vފ���8��EՏ�-�0�*7I˖jI������CRk�ɘ���yB�H.�VD����<��w�j�a�
u�΂��+r��Ӷs��$i��+%���I��|7pϺ�ǹ���x+j�~V��d�����U#���L��/��N�[�d6x�Hn�{ZG�!��e���o�݄u�x�����I"����}u-�j�Q�)R�I���yu<�l8L�A�j�h@ O��l��rb��L��hE��Q��9�MP͍���8d��ޟ��t�|=����5�L��G���,&\v�5A@b��gQac���!���+��Es=^ﲭu�v�-Ȯ�Ky���Ug�O���xW�T���y_O����r: >�8�B-���Jb�&�&�$;�e+�Î�#���e#�,�Y��s��5sh86ق6��կ��<3J��ˇ���a:u|h�����Vz�߇~�������o[�*���\�/i$�H��:��F肿(.As�ٻ]�4No�yU	Hؗ4�	�����0LL�N���讫V��ZB���ON�h�����-h͂K�Z�7P��3��EpWO��L�����}?�j/`i&EO����rȿqv��m.t΁C.�:�W����M�C�q���|�a^jryz�8�}@%���m��#��]Y[S��o��&�=5-����i��(��ꑵA�3�'�E���0�<0�VK0.�:�,> ��wG޽$Q��1wi;z7۸�>b�F�O ��D�ҳ{���(��^|����O-���Ⅸ/�$�A{��a���/���䙁���=�%�nv#��798�cАB�ԭ�{�ݴ0��rD��J0����Q�nӸ�$Z���{�w����Yk
��&�eii��n��T\1��t�M�f<�7CS�~�<MG{	⃋b��<W�a�%�%0ܓW�P�]��ׯ��b��CC��ӊmQn�4�	���_/�zTOl���P������u�R�v	1�۵�O��.������q
S�q�\*hy�>R���M��fs+]E���+2��ܖ�~��g����F�K��wb�̅8�傊��]]i��@���D��9Jm�X���o�Q�~���2��'��%��)�v'"_��h�$�9߶�k��h�Ҭ�	�7?�9Ѐ����%x}+9��1ff��!sX����e���$����u��M�vs8kD�Ď��wԜO���y9������6v�q���C^ʲ�~9��h8$M��=?���`���j�:U���)y��"rF����g\��3�j����;���޿C�a��{����(���^Jg�j���y��OuA�sn��i^�jF��[��`e��5%X@մ�X�I��Dp���{YxY!d2�u����L��.%j�k��\��up���?��$*Yu<�MJ���g�i���68�V|����_��;�"P��B�5w����鍘O���0=��*����(��E�7�I�� q�h�b2��˧��-�zg�¡������f�(�??l�O% �t)I�����+����� ً�x<w�Y3��>�ɓ,����0�ė&z}�N��Z5z���T��.���	{����W8W�JP~[ofaUW�2�Q�k�N/���u�D�s�`�-PbX�l�oj�L݈�
Q�zX4�O���g;s���X���F��0����jd��o8�̔�����Iz�yhأO��H���W:-&h��4,���:�]���j5�ϲ��w6ߵ�3��\��m}�@"�Sc�� ��	�&2_>�.�nI�<��s����S����z�g��p �'�1�aT���F�>y�	mѕ�bnZ\�������eJ�q������J)�/�N�>�����HD��-
E�ރ>��������.�c�)���u�Mlc'Z���ai��Ƕ0�rD�S��S��gڸH2Աm����G���C��pg�G�e��牐��[@Q��RêF�"ટ	O������YY���L�I>�ZJ�'I�JRs`a���,�{`o*ȇ��
�V��j�a>�7e� O`�b���3�n�͔�*�'>�3�����&�>���:�-s�DB��$�r��cY٣z��ܻ#��L��o�ñS�ʬN��qf��P�=�@)ֈ�R[��٢��|E<ILy �t�&.Y6��N�t�+x�k 	m�B��7+-�� ro�o�7���n��WL��u�zW��@�dE�����`��3�܋K��Qtap�~�`#;�9���٫{�������p�`��y<�m�`M{`�:�#0IOcW��*��GHz֐�L��{�,�4P�i��돪�q`��t*�hlr0�YGp��B�P[)���;��+$�"�S#1��*�nR1��ۥ���r�d�v�C�`�Y�y��iIV/�47=zֳHJ�G�!ٝь�ힽCOWj��zFu]?��>Sq͒(�
��8!"��D�w�\��c,T���rL[S���'} !b�a��3���X&CI��<;Ӣ<��q�1O�����P���W�(DlR7b����wb䍻�j��AO')���3eBs䌨C�N$^�)�cm�>xQ�ٸt�k�q@��N}�ψ-� ���0Ug��)�NòN��0?[� �e;W����&�\��\J_,�#N6�	F�Q�V[!�$�$��,D�U�ְ�V\��[0��,�㐂�
��v���с�����L������{��I�a�c��d;�ص��QXI�"qWq�Do'+�,��O3� �+xvSEմ�8L��	���(Ĺ[p%�\�#�Ba�o�s��
�
��V��翥@O��d	����%=(/�^�Y�&�g�8���e�Bdyp [c�Y�`�D���>���a�T�����b���>f �|!2H�|`���Js7G������{:<�Ҡ`~I� z�SO���EZaE��vY�A�X��?����s���h��P-R��"k� �(�{�W�9�q�����?'�mn��Qc7JU�R,*�t�]��Z���Y7�<��Ԁ�T:f���lTB���CS�\�H�%��Xy��-�����ހ~�9�'A6Cd��YU�s�E-34}
�T�9/����d��:�X��t���O�V��N�9�C�M�o0'����.Y����0���z���>���$G��Ƨ�ŭU�aT�4)���,����gX��h픛�pqn���j�9]Q!g�n��Ig�Xw˕Ls&�OE�b�A�sl����V�&��tezb%�7���,�u�?�0;5:C ���	�{U��첎v@!�uR�o��Q��⤊�2(^�����+{̙4D���[�7�X�L��1	TW�.$K�J�H�Zƈ���t����M�qsVAeY�������ؾ�x>�,y��{��T4���|�b	8��}�PY���s';;#�ǆq��S⁂Ww��z�w��t��OI7O���x�z��xc�~8͜Uq:�@T�{�s�ګ�'Dl�h����6]��]$�?��.���]�;�]����?LAg!�*@��2iҦs��g���߯���oI0�����o�R��^B{�zB>,Vd��Ճa�9qFoj��U7I�ܣ>'v�d���E�� ��=\˅Q�`�=�g�Y|�����j����}rƼ� \�$��u�*:�(Q��et`{��GC�e7C������"��@+W08\��e0'�'�T��(�{������Z$�u��X�9*f���f��Pv���&\c�1���7���8(΂��*�5�g1jk"ޜh4�&��0�rL�.���Ro�O��w� ��47���"�Fv���/�9����.K�;�	�y؂D<�ڹ������u�,�ԭ�G��T����(��x�1�<��Q��ϛ+��A�C��̝�UZv�mndak�~d�R�l�����4��Ђɡ������l�'" =a`���.��t�<��V3b�;h"�y�[��n�$Y�ߨA�*�C������S���&�L�=fߛb~p�U����f-P�ͷ(��b�D�׺���!�-�������/�n����Q[�eL����a`ˬ'l�
�mt}�'���3�@�TG�Ka����3J-�.��ج��S��JNP� ��}��}ݘ)�ʗ��/���2{m�I���;�]>$w�>����k������+3ќXVIܟ���&D���oT�Y�sݣ/���=(��*;���(�DO$����b1��������R��\]!� ��ڝ}$���7e��a�F"M��c%Ciw��+o��6���]�
�<ށ��:�lb$jg5d���S����R!@&{!}X�m+u��K�B8W&\�� H6�r�[�eV��
4E��oR�U6W�~�:��u���,��<�_���$���ˤǲY�Ӑ*(������_�Ԭ�P��R{-�H�EiL�|�T��'�#T�EۘF2vipM�>���J�w�W)��m����e�,���$H�Ǔ�ŧ��[��[�JZ/���y�";+���]ݑ_�=[�lb��Ą\S��syDb�s0ƷØ�dI�7Ý����"���q&ٟ�S~?���l���yR�S$���`Xc$-�l��s�'t�w2h ����xf�n̫"Z���~\����֝����7skS���V7Q��i��.w��:e)dg)��WYd�1	_K}$I"Ç,�|�v(�&}w8��s���4dbnE�	�Y���P�2#'�OxwYq�L1�w)�i"Z\��S����
�9yN��]�2��22e����u3����G^G�ŭe��T�v}>�O�G ��O-���O�`x���ї���N� 27[��/�#�AL����k�mh����o  �F�<���9j��`=�Os������3�@�a&�ڣ�a^��-����B�W�\��?�tcW@"	<ÿe�����LQ�pZUP����+P�T+�Ю��!����L�{�I'�t~��b"$���o9�1�D V�+!�+��,��2/5����4�{�4���;�����zuO��C��D�|MF&\T\�4�69��:Z�0eG�J��lv��x�;"�e�'������c�W����Hr�P��Ӗ�&�s�O����BmMEKx4�$��RL-��L��)*�~ B�V��^W�t��䃅W+9p���e7��p���Uh2?)M���Y���k�9?a[w-|�����G�X=7e��m=�X �MC7=����?_(�����~].1�ݝ�f����rƿ����E����V�0��'�7/8º������i�
^�X���Z'̣%�s�U�uy�N�<M�����qR�n4(�JϚ/'��>�T�����2��jj���Y3Z�{D���%͓ )_��ȉ�7]�VJz{�l�����g`�[�L	���&��"Z�K���M���jP󣋻s튮=R�0j�<�V?]/E����T��Fl�'���T��y�BEW^�DѫT]A��U�)�<�.�#	w乖Rk�h�ط���B(#�U��ةa	k�:�@4������FY���-�sK�:Em6Μ
�݌������1�˧6o�2�� 9p��S�K�aD��m�j1���M;@��{��œr����im�+C��^���$���}�=����!/v��h3y�о�-��Iу�M���(�"�,c�𶛕� �*JMі�LDqo�L�iz�K�Yy>�
')��!�_�E��t�"ҁ1Do��)��A��~�x�B=dJ�IJ\]�؀�{h	'�{�h��%��x�/��}�T�z��E�^��]�t�jw���}�=���f7j�2��2����Ԑ��v�N����<�(ӛ��O��c ��F`�g���"�`����Њ�wΐ��� {уf�-��L��ķJj��{��sE+��#�������Sh�1D=�^��'#tZ��-5�8��R��d+C��HH���1r�+�	�ā��BŞ�T��w q.�'��(�ɏ�Lu�,�s��I=_�z_5[�h��:i������,��.�ϲPC�>�V^ b�r}�(U��W6}=J'�i����W���@��n�L��G~��u����/��nNFP�$���W��8�䪺+ҧh߸\WVwǧg�xBE�T	F��� ����������;x!������c��jsk��9��h��T-�R~鼅�#F�~�5�ʏ8܀�����R]0�s�Z�sc�@�����*
E�o��)�L$iWl��YǁD���3dE�9�}��L�����*>r���)�Ӵղ���=�aJ�T
�w= 9�RBCD�v��^�	t��e��7���=�uwY�N�w���KXp���.�;��� l�����c�c'X�\���7t�Z��"ey�����i*�$�i>N2�i0HV�N�`/�n��X���s������-��>�Сu,ߟ�;�M�}��=�z6jc	l ^ q�8~��v�z�wu	�$�T0�A�X2��2�v�ZUzؓ���y	����g��\y��0踺�Μ�|'��}W�|��bv�6�zP8��[�{	nN'˸�7j�)�O>P�Rv�E���kJ;p�='g���W�%^r�k�cO�6]�-��^��ʔ���"7_~�cb����i�~B,������p�dN�[se�z3�}�)��Oc�n����Ez��oB��lG~D`�}g�XoTۆ�R`p��<��u{�a��:9��H A��>��V���S%Ex�q���4���zM�'3�g<�R�[��-�A"
-���o5��녞���|�Zi���1H�9��� ��U{DN5�N7�xCt5�
Vk�����n��(I%-�����r&@���{��y�P|�s�5�.��GQM�iޤ�KhbE*Ǵ
@:;�J�>0��o��-�ƛ��w�ٔ2y8s�>��EGC�Cl�49qnc�����C1��1Jo�����ڄh6[s�?�RG8S�b0o�Qi��bF��ދB�)�C�ܤ��y1n=)!���B�kF�c=�ͱ�j���D!`�5�0, ��@�K)p��.��Vॱ�a-��6y8�螴6V|L�GI���5<S3m�LK9�σI dj4yO�XT���Vk���X�O��P=BIL�@$J�Hx�XlxV65EB    edbc    28d0����J��Ne+����\CY_��OI��	Y��r�\�LOj+�xȏ����M�v͈�#e�q�4�iTf�]��7?Q�Xu��n�>�mha�Z�ZqT�;�3��1��n�(ن�0!�I�틎�a���X��{u��ؚ��b|�ĹlxV�;l<)<��������hF�.�ɨ"V���_[4(�s� qJ��o���vΆxroO�lP���P)s�������6_3�B�WK����%��\������������f��B9�x���I�TA#�M8kz��a��S��j��}^Oґ��XʴTQ�ȫ�т�1!+֚g���֭���-w���rN����L����6(őG��69��J�A�^��&�dojɚ1?�g��Ⱥ�Sf��2v��K��Ò�����o�5����&`v��ւ�jH�e|iX���$�6��Y"����X��5��S.h��V�V�2B�����\�Jץ/X_���k�D���-),0)q>$�.� �]h��<�\���>9Oz�l�'����t������'j��zh��3.I��ew�Kr��������=����Ĵ��uį{�<�U�.o����>P��(�_MO�6�=r�ώ��B������׷C�23:�X�˞ 9<C��|���F�,ݍ�	��ՅUHpjG5A�������h���!	z����J+Xo�EB2�0Q"�D��b*�yTvgR���Rg��]9g��ɯ�,��#5F1�=���y �F]���gb<���iy��%�4Y�@*�ܑ��%˴��#��R�u���_FH�b��D�a����x ֚W��+�q�G��J�}����kU�+�g Wё���;4�¦�+��J4d��p�ĭ��5d �����2\M�Ǹ��s��x<]rHzN쒥+�UO�r�B�YLpq��U�J���8,�����X �	�z�4<<�I�Kp�� �6^~s6f��������+//��|s�!�0\���c? ��[���h�?Y�6(Z��`p����2�����J�٩2|1��J�k����_kۤ| �OB8t��(��Wy��m�Y�\�_��ZB:�ж�'�U$��U�����KsN��",����Y�n����.i��Ӗ�$>r����~��אi����J+�����re}Z��0�er*��y  6�4���iwփ�>!c������q.����\K��yC���(��u��Jv�5%))�C���v2j�sڋ="��c��$��牁���I4z�������M�&��I&S�7awX��������6^�P���n`��T����|\'$�U�E�@��nk�L�
?�V%h��cA�M�[�����vC��6k۰��s��&e֩(ܰ�V���� r,y0ǂTc9/�Ȇ�B
���h����:Ӳ1�V�?�_��&�S�J�h�~c㮢jKy��ӁGV�]���k��LF��#-�ۄ�.	sg����:��`ULI~L���"n=Ԁ�e����r��_�o^���k?k����A����	��֡�g��~�����[Eaľs���h�}��̢hO���Ƌ�	��ݾ>m+�S���EgB3,���W,BC��տ�xȺ1�{�,eIw��C���O���~�ƕ�s���y���|�A�s�.��,�s07�c+E,��mS���^Rx�өO��A�w�D�8�`1.�=1��!P�ə�5��Z3r��4��
�}͑�)bO|FA֘''�;F�7K��<���E�+`LQ����p�H�ؼ������a%��C��1" M�����dm���VL�z!mOmSE/���c�����%�s 垨�v(Ɵ-�炸��1�f�@Ɠo.�5����&�+�1�N��Lu�G��عS1����Fɐ8^�g��3�FGt�P���U&�a��׊�qb ��'� r��E���$�����w;4��u�����D�d<�x��߄i�b��ZC�0�+�~���F&^ETt4�\�Rf��jt���Մ��D`Q�0���b {f���c*Ƞ�E�х<<�X�J!8	���'�<�����y�>^��x��!��YL*yS��;$��Cao5P]�(�RDQ�ࢃY[�]t����#�HԐ�^v��uZN%��uK���0x���&�J�`֛I��d'c����.ȏ!]Y�i/�_��M�S}g����`��_Z�.����ϣo�`�k*�:j�b
](��ZZ4�� x���w"�M�jG�[ 2ۅ.�X�V�#}߁�
�EM�9�nb���
�]��9�_��!��#ە�LL$'>����ϋɯ��(�!�W��7<��X�/�D�9l�n��1�d�+�31���*�������� <��ӥk�&��R~i� �x6<�V�������\�������?}�]䈏2�p�Ѱa�)M6��Da��������QT��I��>����AfK����	�e/X�m�mI
]�s���~\u�6=�Śc3T�Yb`��m�|�M�8����M��'��SH-S��CxN���.�k��>�+���2���=`K�D4Z3>�"�D�/0+&���Q|M�}�׺�z�=���Zދ;��g�����vU����P����h�b�xvP�JY�ɱ�"3{����&Be��C�XR%<�*�\�014k��r-�N��Z��K�Ϋ6����|Re���.�t6��3ɒ�T7��%}��ihP6_]=�s1�����C!yG�^��uŗ��K�z�?��3+��D�'�|��0&:w�8�����a��oVXHl5�GK��MQ1v�t�qz�sE�ZIK�W�u4�H�h1Ta�YK�N��f�fޠ/����a:��I��Y�q(���t{���;�3P�CS��f<f�L�ޚ��O'�CV�jt��b��F�PĴ�M�XO1���
q{����C
�g�>'����n�V�.#���	J�HL��b��2Y��.�s$1r�c�+%��+�¯�pYv�G_�S�k��&I�߸�U]�����|5�
���2�Lj_:�/*�-c>�X�t�YЈŝk�����n?:.p G	ߦe}$ms�c$Hs#�^�ϡ'O��y��
J^��)��o�^�|c��]�#�Ee,l4� ��<�@�]��e?pi��t��E�?K !o&Iz6�m·MI\-�$���+WsUnܪ����X��&[3���_�,cp��V�ƭ2s��iY�$B�����gD�7Ɗ=0!�AC�@��"�]�0�e�}�ϖ�����-l3~�k���q��Ġ1?Րf#z�R��.B��H~�s�`Hh��K��ҷT�5&q�g�!�.�.���@	���P|v\d�� V� <�`�>B��n��i;�h7�_M���k)c֓4M�IQ�N
Gt�'�6rF0�כ�)�8v9�{�o��y���O5V�u��;�9�ټA��*�" žf9h�J��v�+��g�Zx �]�S� ~O�� ��,�����8�hlJ��,?`���_KR��z�#�Kr���k�z��}��2H�<ۗ�Z�=���R���|0�?�Z�C"����Zs�$��?���Y�X3�'px-D�y��/��-zGp�\]�H��D���@��ҝn���)j�/�-��w���n ���^ča"�l#R�(^���[��L��q��ߘ���OlE%��X�RqL����R��2cL���Mᐻ�����ܯ����/.u�p����JNa��C��*$4Y���\��}��5g2f&���G�����.p�N&bx�l+O >��ɻ�؀٭�Y� �u?cz*3E�s�G�1�4�z��f��=��&�6�"�XB� vw+�D���Yy�] `���[H��fj��VL�:��+B*�V�i��U�c�
�b�/�p����H�i�tQ<�s5i�G��:�^c>7�B�V�	��9M��ǢQ@`�.�b�zS֥�3�ϸ��u�	��:7BG��=�-�Fg �p5���.m���~�(f�����q"�uF4XǨ�k7j�*T>�Pt�a�K�F�+��-׻y.�tJs-�j�T�����b���l�n�[�H�g7����j9��3E�Y<ɛQeE>M�6��OW"!ᨿþ���͑�)y�x�mC&�<����şNR����H�<8\L�4�$[�ͮ�ο��D�E NxJ�����E)􀈈P��?`%��#���z��;w�?Ʃ����it3���E��Iy7�*}�M�Ӌ<�	M��i5�m��D��������ףУ�0�W0C2Z�{VH]����H���՟�E/ӣ��L�NO��)�h����}^}7<�'��F�+N<zl���a��kN�8��6F�+��-�'ǫ% |O<�e][S��=}Ri����}Ek�$<���;UE��o�i2o��E�]���l�I�Ē��"F���2̌Tj��i��1�����$�˙�U:w��r�����q�{-f�5�¯�禔/�|7=��t��P9.�0���fPU��˧1O�1]��6F&0���;���]l`R��̷|�
�5�/K&E��AɁ�c��ۉ�a��x����C�\�06���3s�f�_�����z�Cޑ�}�s�$.UZ�'������	S�0��|[:(��3�r��i�����?=�$#��p �P�!!V��`ϖv�T^c�֥���}�<�c|�AG,��R�0��B��^5�n7l~�L��#hë����~'P�[��e+$��;��@�ؗ�-���ܤ&���յ�Y�&���A��A��azۑ������GЈcry!�L/�mW�1����6X�i�l�<ʺ�J�ț�� U|����%�w�qsN�My/����>"��zn��]��j0[Ǥt#U4ua
�t���&K'"I	7���1T�Ymo6G��~c�y���r��F�<����V��پ}�2�T�G�.��)n.�k6	�;0�q`�3� I^�=�#�og�~��� ����~�Mq�&K���nTv�\����\��%UY����1- 05��2�J�lB}�i!3�F��cܱ��q��西��V�,��6ޮ���zr����	����B���
�qa��5+�6�G:�m�S<�6�v�w��-R�]F�K��:�3���}�ǝ���iE�C΁sCx@�u]��C>�e]霭(oҢO��V4�Fѐ���W�.���O��Q��L37���>h�]St�9���	d~��W��VZ�y��f��@ܼ�m��$��G#���R�Q��;���P�qjx�I&���8c�3.ܣ�o7T�{M�AxӲ]	��B-�X<���SQ��7�fl���M�X8��̙��8CO6nT]�;�Wt2y~f!c��(s��oR f��5=:pBS�|@�3y��|������  D�����V�]�@�aV'���C(�Ct��X>�!����%,)��G��Ľ�ab���� 1��%9�%+�����F^͠~�H���6@�S�1�9������Dw����:?`��DT�:7��|D_��i�Ћtۍ�PFRAT�8͋-K�:V��3�h&��� <;FZ��-+��j�r��G-'��w��'�ۻ�@s$>:A๨�W���2�Y_�Y���	X?SZ��n��*rC���1�G��n�a�g��Iu�$K�sQ�z�Os�y�p� `����Ztv����hcf�M��ґ�N�:F�;rj�d�b���:5ҭ���,���:X�f�@g���H�:T��p�}�д�'���%_l��1W���U�U��E+�������)q��4���6�������Cp5�vg���1�P���uο"��[4K��/7{����GM�i1:*�G��z	�:!�KZ1'I5��S��a��zi��� ���M������x?�ТU��&���yf�f��[ ��Z��u�S}x�N.>�3��5�uV	F���I��ls����E���������j��$�^%"��F�?���nZ�*!�zv_�% ��Ϝx��?�s�$��(�|�S���>FZ�� ��)�9�UtvM��F��˪5��EI����RQ&v3VYOX�tZ��U_n���+�����)Z:�>��e��c�^4h��,���ᔠ��`��y�c�#�����}�����o�!�s�H8�ɘ�IX'p�8*�^������<y�5(�yM������<�D:v.���|�	���Ak�+Ɇ���iW
�x�V�0�QSzn]t��J�-R��-�ܗ]�����%X�4�&*_�t��Z�%�g�SYEJ#Q�����f�4�M�Ir�qV�D�sc�aR�]}�A�%	9�K{4nQ@%ps ݭ+���^=)��z��	H�X�"_��	����C��w�]�^~�ǺO�U_V�"���a\*X8��{���Wá��L'��C[!��1�K�����.����8�	�l۟4�&�YiM
v$��.��E5(��?��9ǯ�.<�l����_|�c��㨌����mv�҇e��z���40�U�0���!B�o�F���Y	O�[�~tj���	6�@3)�ot���Z�m�9�6�٤�9 �vup�3�����±:~��'��Ά.���yG����>�Js@߬����,�T3���������a�l��Șn�Y��4B|%`�Gөib��iY(��q������$�� �S. �#��KC�CzZ��J���9�p"G���yɌwg6"PB7 ���g��Ɉ����z��V�I��$�)��Ȣ�ɴ��,w�3iӒ����j�2Жr�`�b�i� d�O�x�����1X�K��g��?���B1�P�بF�3t���$t���z;#o�U!$X�����2����L���w"лA@��gjrC�%W�� ����{�Cw�
�8f�X��vw�hl�k��"�b_�$�.�����?��A��BfQ�JV�`�o�L���}p�������6��7N��NvU�<T˚����?=��ٙ'6o|Ի�]p���ڝZ�cZ<b��5�4���#�v�Ӵ�ُ���~���T��un��$@�׋���p����\U�wŻ��wL��}b�Vh�0y��y��&����VU!��h�B6.c�]]e��T,h��4����O�ƊpD`Ī���^|c�;gK��@��s������:����D����+g��V�B���vYG��+r*4\��%�RE�ފ@&TQV�� ���'��2r�hB���$C�����X�e�������=�����m�W$�:���r�*�t]���R�Zޥ؅ͪ+L�$Vж���&8���������{���o�N'��l��G��G���~$�>P:�H�M�ͱ�#��ˁr�r�^O������duz+��:Z)7��\��@�����L���>|���g���IL�^
N��,䅚�<*B�e㹎���2M�@�P1'D��o�2�J�oO�� x~=��]4�V���"�D��<^唼J�� W"�=�l޸�XV�י�h`�ha��(mOׄ�s�˜\ҦQ��Zԋ��2g p�"�h��1�`ɟ�WVq����t
R�.��%Urx:�Trޅ��~|J�\���Ä�:+��Ct{���+��:���{��CM)�Ê�R�	Ҟ��wb����.�?�u^�'�<��������c% �HǬ�R��y ̃�Y�	�H�n�ur�L`@24�Q�!�t;iK}x�Jn���C#��ϒ�&�Ð�V�-x�]�h�68/_(4(�ܝ���✫�p�1�WQh�Cd�Z�[zr���ɘiJTD��6߮lb�qXM�e9ǃy�2�Q=-�U�aæ=/��(�;�r9,1:?Qs:Y-�`�����%�J���{����]�~���X5���q
P�}|A��p����?fh)Zo���>�[�[5��6�0�y�&LH㶝YY�;q[�bV�!g��(�m�R����)��x�xӞ"��=tï�`������A؉��
�.9� ���{�������C�M�.���D��oh�$֣�}ؽjc]f�����|m^Ţ]=��!{�6����g��9�#k�!��-[��4��fI4)�g�0y�д��o�~`��g�W�B�wk��UD
&S�p5���7���Z ��2ӑ_rן)��y����M����o:�8�ހ������!�9S.��=.��Y�p�gFW��GV�<0S!ZZ�������_�F~pJ	:���<�U��Ŝ�sKD�.=�?
.5����6��ǀHa-E�.d̗�F;�+BK�'��ߚ *8� ��.�,I/��� O7��}G<��ٗ�K&X��׿��Y���-~S��Sa�R.Wf��<��s#&Ż�۞4�-������G�K�GU��ҷ����5_�x�]:�Ilƽ(��!
ܕ��j�ԫ��oa��,�u|W6��ʡ�s6on#���5#��
(~����83|��V�aj�q|��ic:%��		A��2���������tav��j/����<57�;'}C�"��2�H�\�X8B̛���F�����h<$����vloa�,4��mz�5�+Nc��'E4���3��~[�LnN8]`Ft�\q�;{�P�NJ��9ٕfa\ϕ>�'��m�AK�L�1Y�W'{'�� D`9Dp���ʩ29��k�y��s�=ī��1fc	�����w����x[f�!\JDJ������ցT'��.ӓ*_�vK�$H��2�n/��NM,��Z�=�J9��LA����v!~��Me�\f�HPwX���V=�PF46>_�����S)���Cx9t�	�i[@AҬdd'%�v�=Mz���5Qe:!2SKN|����I�����t�&�FL۱F�����C*���׽R!;-�_��,�}=��i���SI�?�NZB�)CHo�v�3�G�ۊ!��?�����Vƶh�������=%�!D��U<�ߥg�=FEɎ�e`���c%�s��݇\���n���6H_.�Yq<�롘�5���FSC�	���`D�?W�3Fn��i6 4��O�t�U|WmlS���v�ga"n4�&&�.�k@u�ξ;
X�(JCr�=��3�!���f�����-W� b'j����X�}��P���R�Ƀ���=z�ai>C��\y�PV\�:OX��� �uKe,�hi"�����z���'�(\�[*�\�pS=�����_�ڪF}�'�����Q���&fq�ь���JA�ğ�d� �n����3L�{mh���h�+hFG��<��~�r���{��ɴH���2j���/{��u.��v��j�S��چy��)ⲒyV^��+��vq��,�3����\����>Qm����6����r	r���߻�av���u��;Eb��û�Qr'e�X�rF���v#��	����}U�w�{���{�u�QMwZ�u�c�-�ǅ��v �m�����'��C9r�ҧ��
) ��/K��� TLK��W�o$=�r���*i�V��j�A�0��p�����y�ӟ�	�p���PqiI(կ����pr���y���rZ;ie���:�T/H��Ih�M�=�ߜb�~�-7�FֺN�
����3��5������У��s���(��*6�|��Ŕu+@Ǵ�ŚUGސ9�4�҂��P�j�$f�YV�O���(�E<�Jֵ*��+�x���)�]����=V��L�3�a�����Ǡ��x��RJ}׭��)=�t�
Yy�I!)J�o5F��52<3��B�gȀ�z)�����KS�䬐��OU}0�B��
���H	�$���8՝�	-vs��?jfD�:s.�>���f-��;yb�V�Hfw|��ˇ���z`�������f��N�� �F2������� 9��.�|>�����Y�/����ɬ�&��0��~$/�sB���x�&�hY���e	 Hxq���F+�%��/I�bJDL��
�q�;��܈q����e��Br����v/4����6�-0�Iٓ����G��b��)@�1/D�7�	 4��[H��/Gm��|}��Md��i�BQ�7ʖ֌���/�V�����W'��ѐz4_���i��l��A�A�L+}�[|�NPv)lǬϕn5V�%��i��e�2��;��i�+ui�\�"����AD�����9>BW�ݥF*���'%_}?D���H��H�tm��G-0��WK�@y���S��
����SW��}\$��n�u��V04�H<�S�M
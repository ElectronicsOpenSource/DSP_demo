XlxV65EB    fa00    2e70�a{��Z	�Z$���T3,����!��{�#3ne7=���X�{������X]�2��8)�����	���(�\�,v�L�v��^%����d������\\W?L1k$w0Sjo�#�騢��������w`އ��n��	�ָ��'�#�Hn5�o�1k�z8c�����
������0ge�����y�6~���r����`�b� ���<f�N� �1�h���h�2������%��[��f�Kd��)[.��C\b-9Cx;RG���a~i�Q�h���&2���]f3$�p�h��T_�zJ���#ӭ*R��a���>*�(�ɏLK��ah�yT4s��ݫLF�A9�2Ce�<˃0P$���jU�*+j�7�����^��Xr���E�=Wjt(�NZ���`DE����٥^�4��O[�F�y��D��~�YE�%���,�6��
#�I-ވ�;t����k����5��uw��OW?���(�>�R����Dt�h�|C�QJtQd�9���E�J����4��Q�������Z%L�%��f#��1î�y,a���3B����JP(�	;���2ı^9�/�a
��
�G��u��߅`�Y�mIY��/�uPqo}�]q2���E�\q���|�f��ޛ�`�B��iD���1bH�ۤtN�a3��U�Ouk>�eXw�<C��e��������N�#�;��#��k��g��y�Ҩ��v�i�+��N~x�w�m�a��N�q8Tb��"Qㅤk�$��t}̶��$21iJ""��݉IQڌ�9@T�ge��u�c�w��X�oNi�"Q�����zN,M5P� �y�v;��!kyp�'r���;=�UEY]Q�$�`��,�{�g_
>��W>�ӹ�4��&��R�+��e��Ol;QG���Íx��.�Ǎ��W���-B�ҡ9ݡ�L�^'�f
�H�Tt��HD�y�JP��A�XY��� .Ҭ�(B�d>w�Q��qm�qV����]1�2Ė1������f��@8M�a��3/SΔ�S#�N�眹��|�V���?�˲z���@�>���x�
Q�b"��-�v~;�w'�SԚa��0��z�C^=�!)n�+ɒ:�j(�q�h0D�6�A��1�N���<�rҪ���¯c�J�X�X((�)�CJ4WnM�z�r7W:���"����\��� <b��ᖪ�ԡ yh�Z���d�7����������	fYbI8���]��֤t'ԣ�맹�i��N�<��`��!7ԝ���=C�l�,A�a�Y�ж��Gδs|U��w�K!I��N����/��<|q�eu�˂�ސ��1|*��t������nOV-���2����ARy��=Ļ��o��������d�M��ގ�N.db�da�N���$�E��1���\Ы��a����Y�&�R����O��RD���΀�r�"����z����,uj���	!4� M,�����A���:.�Z3� u\!�UM�DŨ����u�j9<1[��1=�h���Δ��?�����l/Pl��ϕ���'��=��ft�����"%���I�`��C"
��!��j��@��b�n�����|�e����meM�:N�?�	����ͻ�-��[2'�_�'AU��(���#E#W�9�~C��|�X1�5���
�� O��3���/�䷔�5�Z�Gӊ۲�>�:�_�.N')`�9<�!���<�k��k���MM����/�?�g���Bϵ�si�Qzm�upF�pQ��h�\"{o$�����t�Z����a3rF���10Gn&󋠑�xb�?��X���9K0b ��d�� �ɶ��*�$�/���y��[��������hD*́"��`-U~�_��0U:7��1F�rt6�5�B�����(��t���+?��7��@e�{]~ф,�g��~�ْ,�,��F�.���&�!���i�EVƇ��GY+����f�OJ��7���z�ΫN��̀�����ˇ��g௰r �Z����
#J,��6��8�$k"[D-����zH���;v�wQ�s@/(��L���+���I���劧�ӑ8Bo�p W"ϾS%/)�garV{3f�4������"D��/ɏ�hA×�dv��͓c�(źzS�ל�cg��L��?���-]\x&G��;���|�l��He���q>z�Q>"j@tQޣ��$�j���#���ʕW���&bJXnF��{O���C}TVA���R'�C������0z����xD���U��N�C��zU��,�T?�e���wk�f���<~����N��%���\�\���,:�P�1;�D9t��t�f��	���Q&S����q�F�l^o=��7��aY��`���1���G�'���BM{A��r4O5j���-��K���]y�W�Q�m��U�5���?9�X)Q�����Թࢭ"s9���AK�p��ޘ�6�hi�րU��([���6H�B�2���b�ɌUਠw
č�7�YGG>��b�C{Xx�0������P��@��b�'gR ���arZ���f�nu�p����tK
�q��R�u1�A>���~����]�1�!$|���U�d�&`��rt����#$ӀW�0[ٟ���������8m�P��^�
�mV	�������P���2Gt����L�����r,#�І ��YW�VewP��Dm1<�חo\�\$��;T��e����L�]�1���]������R��~ua7D��}��X�M��'�s�S��/j�%�Y��؃D�%�i2`�w?���cC��z�����;^�Id���m�8��Gr_y��z|acR�ᱪO,*�V�'@��+�O�f<�X+%2O��71�f󀚄��e�r��9b��"X�|�ܪ-�:���9���B*R��^�.'�t)
[>�T�Oc�F0a�{�f���f�ڱ��~����O{t͍���h��l"�ՠۧuEY��U,a$�%ECt���?�9Q�!λ�5����� �f�plY%arϕ��o��Y0����R�@�Q�f�枮�$�
���d�j�QO)���g2���T���ԟ`��p����ʷ���e	w�*�H�e�����jAf��A6,	>A��ň�W�&��B!I��.ʱ�����Mk P�S�����ˇ�P٥y�`e0�0�bv(���t��~�q��w���D���������LT:�;�M>�[t�W"h5���2@��ګ)���
�9z���̭�21���~&�Xq&�wVR��]Y��0�Ș����s0ѿ��J��" Q��q���'�L^5S5�5�+0�����1n:�8�������O�����P�%=hqA�_�Ͽ���ʄ�zʛ�	�wW����V��=Kyh�.�}��;���j�n�Kx*�G  �  � :���m'��	���H�<��ۇ�.=F`i'��U�p|2~�`�����:ʟ���^qlH�=2{Ox�MA::�������i�y�_"���5'M(�X�;FZ)ku��z����͊�j �
�8��4��A<X��A����'�P��$�TS��&Px��%�+�Z<~��|Y	���M~�g��<_?�1\��	����_�����NQ���ܯ@mKc��ǁ��&��8Ы$�wQ��d������DS1rU(��r�C���|g��~RS�j�B����x73:�q`�I�B�=&�yˆ%����K�y�M�*ZE�ODFgk�Q���i�)m�W�˃~s\3��"3�7�=<��\d"΅��|��>�m�o��$x��RII��w�w<b!`^'޳�<��<C��00C
�.���������/������
6�T@v�<^2���f�$�/t����X�1��n$>3Q�og��Go��h�璼�Q$zj�3��?9��]��bٹ�sY�j^�<(8���?Sr�.�[��z1�k��*�ʣ��럸`�$+g��T
�����69Gy�QmE���J"��DLގ�_��h��Ҵ.��� o��Ύ�h~�Juʢ������|�Ps��q��bV���;G��QZ��~o�`'� K��<Z�R�@������<?3�7aA �/�k���K�\Bg��CM�m����%J�h	��f���@�_����%��~t�ڞ)n�_�_��f�s��Z.Z&���-�Fix�a�ՙ{�c�в���u�P�xZ!s��ԕH��'�~g�G٨mՃYj��=+!�=��W���t й�(�4��UQ�<���;���)6멮�±k?�5��L%fp3\c���ÈMյ���;�l����W��>�XG� ��Rݶ�QR�5��@s-h̘� ��`k��q[��(��W�R)ᵡ'��>wvF��KQ���UPn!����ɶ��n\U5�ú>��R�R6N�aHY8	���Ks8�g�+cUI���ȭŔ?����3>qa�>y���y���t;�������g����_�S����_��u�w�:�7)	>�	�ֳ�L0�I"1-�s�}d����*�lB�l�w���%��*o@�|�`�� x�lɔ2T��cL�)J������g�m�
 �����(>��*��~U��4���� �L ���pG�k1n�5[A��]^p�iT�)���C�&�7=#��Z��g�~�?���=�;��;O6�6Ɛ�X��F��@��w�X�� �J��Ӆ�|�{�mN!�cFF�a-U�w�I�r�?�P2c��k��3D�b�9#>$w=@�+��=%�LE�J�̓��7��ӎ�}��Y�,���MF�sؠj>� ��Z���\�i]�8��Dr�(1�*5�-�K�;�B�1����n�Px�;����^Z��$��>������Y�t���c�q	]�YW�1&���>����u��^9�Ҍ۞rH�f�s���P��1��ّ������of��(��U�n��p�Q��)��GT��㦿X׎	?s����Kϡ^��P���Y6[&�ydb4~�v��>|�-��E�͖R_j
x�3!Lfp�5�(K��MvP�1!H�x�1�)3����E�{9�8���}�]������e-|$�ݠ)�	���iܴZ7��/b�Z� �'��/�5��#i�|S��/�l����HU��a���2�F#s8��p�;{r�[�/T�;*��br��`��M@�.�W� %ɟ���)��a��mL/��Ƒ�Mp�.!q�5}Z7<C�Tu�>v��:�j�Wve ��T+I��T1�jv���+�����I����ݘӯ�N`Tu�I�0���"�<B�s��4^�}\	�Z�;��#�zc�N��4��k��F��������I�"м��wvZwN�~&ЮF��@2�y����J�jw .;����s��`�I���y
s�QJ��=��R�|�u�݊<4�� ��>��dx�3�o	��s%�j�&���"�W[����z%rP��/���Y��[k�%G���]���r�.X�x[��ԩ�r�J��{�`b[a���uvm�%-+���q��4�ˀ�����f'������U�kO�S��D�`�L,�0��5A�6�C������@H�fJ�۵z�`$m&��9M�7��x�~/r���.��l +՘5��}Z�	���IFo�������0ji�	��[�;�0* l����>t���_G]n������3lZe�d���^9����Ձ�>8h���'0fmnTk� �f�V�R������v��@��<}��8�dG��g�C�nN��h)�ī�K�`j�'SZER���0����UC�H�讳a"L���%¹�{�aCÇ��$��h��u`����:Y��~��J)��`{%�9�V�����Y$+)0us�q���m�h���e�z����j����C��]����r���'��Z�jCTj��(��#�un:,읍�Nm���}�HvS@{/YHO	+`����0�:ٽ�BU�J E����,r�Dw�,R�c�n!CA]��^��\e� �G(��^
�c�[��_��ȳ��l�	�)�������(���߇𱗩f�Qm�?����M��v͗�M6�i���p�D'S����g.� �g�vҚ0)�[���/w$�_-��E����yn�}�4��j�F(����se�E�/9�^�֨���G�j m��vB��	�һ)��,D��T��9z�!������l?����I*�N�#����*v������l�(��~�,Σ^Gt�|8u�:�MDs��#o��9L�XB7����ƽ�[��%jp1-��Vڝ?���,U��*�r�Xi�=8ŭ>V�	g�9�C��z)`:u��\QS�B'��o���Y���&��b�  ni�l��zu��3�u��DUT>��{я�c�~��<U|��.�t3�)��/�{g��+�I�adF��\5: �FG��ʎMQ��DR�Wo%�w�%q%�@=r��׾$:'����g��'�2M7�����l��b�C�O��ث�B�>�̩�i�[%m�1�Y��9�-�į�=�|;����rSt�a��S=�u �$Ȅ�ὅ)��� ޸��դ���q�-�h�g�Ш�*�e���y�+��ߋ.�
x���
�龄e�u�:Ļ����4��tz(*_�{�R.�`>&V�<��)�Ai�[9	`I�۶&_p�ƍ�O����N1���:.���c'����v��X7p�e��|���r�WZt�5�6`D�Kke���(+p�������*Y��] �ݿ�$f��i�l�Я�e�r��FN�k,QD�i���X�I�Sˡ�����oWd��g̱�<:�����^�^��n�J.����9e�f�L`u�`��H�iA��9���A�|�:���Ax qc��$��N�P�蟺�?U�Pu"��fN�J�I(�- і����
�Ac�9��Zx������~�/R�8��k#�Ï�r���Y�xzd�>�N��{H�R94�0+tI�	�e4�ڊR^˳��y76\������X��n>裙J=(�1A�����a���7�ܵ4��n��+�e����wݞH������bңN���z�zLtC�"@Lz��`"y�����<~��I>�S�܃���(DA��<-�m=ӵ�	��t�|ZR���(�,/'Ӳ$���������L{A�Zf�O{!j�WQ�6����r7�X����M-)��^#�č�JY�5��!xN��ע�N���A����6�p����wVwp��ax��5�\�iWՏ�	�Ф6/X�|K}�� I�T|n|�M��I�d����ls�T�/�\�{p��M�1|=c?ݻ�p4���4	n.��~;�K�/�_cx@h	��^�FB&.v���=��\E���k�Έ4��o�z_�6��O�yR�X��_[h�y�M/rX	erb�~vr��UEDI�fxsk~�K�oRÀ�~r$p��*�������6��
�̞q"|­����#h�����:f�:���:Px�`��|�]���&�Ǵj�q�������ϻ
!+ $?1yt�y'�F�Q���u,6�r��~�OS87���R6�����"��L���=�p�I
��P�Kb��=��R[�B}!�c�c΁�������n�?�m�����5V_��������r�"�ut��Cd��n���ύw}�ƍ��D�0B��"�y����/}�p��D���^4UD�ep����<��r ��y밹A0���o@�7��^Ż�Չ�U�j�>�!�+�[�l��Ùu��a"�7yt��i��ͼ�&����8d���"o0�n�0E�B�hK��m@Dq�aYd���v�<��ؐɦ�Oz��]����q����s������U�8٥�%��%�~�����56�+/�dz�c���
5�Z�"��i�=��hP�ºɇϓ�g��"�I�d]:��F��v�.�6�1�:������7/�:����Q�̓�QG�EN�E���#�l�[�%��6�ҡk�<,�M!�|�KGDaW���:�K��yp%$&)��m$����@�*(����ͪ^�3,ꡚ@|T�����eB��E��7�d�ER+��У���[&��y���/��%�g(��ҏ'g~1��ש�D倌?�[���S0$Hp^�N��=��Iz��2�����v�+a�!�
+]�7�q��C(TK>}AϹ-�C�}���=M��7�#�}�
�X��7���G�!�Muc�꩓�oD;z�<Z�:D쳜�%�U&[��cE��s�V*��G�W�SB;ؙH���k��Y�D,ӕ�\�B~�S��v�M�Nt�^�)�0����p�5��ba���|(�p��������4�~���:���e������C�9쟹=�m�5��1`=6�Gy�f�HE�g��ȭŤ�ޣ]�sw���9<c��܎�3Bſ��{4|�^ّJ�lo����P��9��4�/4j�K�
0�D�]���2`�~���*�ax7��H�qF@�_#Fp���c��A��)Vu^20��e�����Q>��9�7묄������Ɨz���@� )E��Nt<�)�)����4��ŖB֥���!�f�c<��]E�0b=��s���'���M���2쎨�=�KyOs�|
lg����"&&�&Uos��	v�A�TcF��biu���B�`A����-�*�ͽs�q��->7�A�$�t��=�;a��z�w�SY����@��;�m���j:�����eMa����ƈ��8�tv��[X��e��b�F%]ΞFx���t��eC��yv/����s���x���o	�8"ۅ�1�%:�9Lj5LYGKK�i��~����ʂ���R!����uN�_M�����-�*R���@����N[h@6CϼZl�Ki�x�q����̮�0��9�b��i��������<Jx;�3��~�����V}�`�y}S�)�خ��H�N����	>^��f�Sٝ�Pm&� �8Uȇ����I��� 3إM�o���ܠ�6:������j�m��{,ٝd�{K�[l;����L��,�E��S�f��̚�/2A�.d6W��Kn;9���y����?���]���0�(;�(kr�V���0p.�"�L�W�]����&�"y�R��CU��:����ܽ���pTB�����8Z�Z9� ��R�XE[|�Xm�V	
�4�*�Ђ�!ᮖ9��o�����A��"Ж&pY�vM~o��?��A£�f!V��~?���
��c�J�9n�~���]�쟂翜��N�3��B�s.$Q�Vp{��a`�>���,o:[���3K�M��� �܈����(�{�<Q��Ƨ���R��2������t`�\<���O���E�[V^�a�]w���#y��Ɍ�t_�X~�-~�jB�C��Y�C��O�?b��t6�F+�h�$��F�����h�i��r�ΛF�1̅��ª�Am�8�-.j3�����d�۟-�y(�R��I5`��c�z��M��ӛ���f������4Ѩm�kuwA�����۰%ύ�px
���j�H`45�	3P�5�������������"��B�\��{e��0�̽���g~������idy.t506d�e�Lp�+������=�J.̤�춣F���W=Z�d�����3����@��J��6S�L2�z9� ����I��4����dl�\���q�i'7����wŰF��Y*��x����z��,pa�G~Ccs������J��R~5%'D�n�5�u�^�&=A���l�$϶����a.��l��P�)̢����c����%A�}�W޿�'�h��ƅ'���y�O#�z4�-aְ֋u4�I�,��w��ٰ���"m�'Zgq���m��|�0���X�mz��L����Ț�KD���/��W�b���nX�%"~�Xvv,^��-��cx�S=��%u���:y�|7Yʯac�� ?��e���je�}�P�<���~��-�*(�^Tl����[;%�Q��X�Z�N�������Ĉ���U�@�jd�%�0�j6�1��uZD���V����e��ѷ���'�öx�/�����f�&�o=�*��3~��D�O�Fp~���7H�q��������R����O60LY����K�L����).��qM�UK�wC�=%ߺ%D��4gl�-�ƛ���*4=�f���C&T��`-I�JҀ<�gMB�J�H;e��(�~�!:Xel��dW�m7%�=T�QD�^߆\����lD����8�pzrHoJ_�������~n�x��}x)֧	��5�$��5� ��ٶ�(X�R��{�vܯ&�|\���L����_i֢�]u���ˀ��ik0�w��2�>kSuq8s/wѨz�4`��i8����G➌)˚� X�)XZ�\�����c���m?d�Jk������*�[�@�i|�zr���m�Z[L��OG�O��){{d,�g&�ԗ��R�=��I#Ρ�V�`F�y����RL��F=�\^3
� WN2-�����ӡW?Q@/N��c�����q�T0���!a�=ntA���I����:������4)s\�����v��P�0��0x�%f�_�q��I�̲�0ڟ����mm7w��]ֆ��ו搧�|wRuh�Fw��;?EH�Jۤ�1�
 ǭ��>qk��*TX8�o�c$�s��.�Cf��	J�T�ȝ��^�w��^����XL���7P�&���5�|?�0�*XV�v�<��$�x�������BӢb�-���R���\Ӯ.��Rܘs9�HmR�!r�)i\��P*�IZ"u��/���	L�w����5�w��FL��+B�P��S'~i;�}q;C��m<�ħ\XD��m��m��M'F?�׾S��ɇÙ�i
�p��G'�_�HmT����gJf�(��yL2�-x5��m�J���xzO�ծ'V�>&�(�(�f�5����I��TGY/v��a�5s`�:X��S���'E%�����g���bT ����8����	��eҙ�]�Һ����z	���10r$�%D��/�:ؤ�Ag.�F����PNM�����ܱ��?�:��HI68��`���C|͢7,�-�s���B)��=o{6�Σ��Ym�rL���s*ɵP+��LI�ΠmK}��/�9�}�z�s#)�������2�bH�$˰N�h����9h5�t:�<�@�6|�u\�P3� Z� Gk���O��>y{�Kеm�Ffn)����jV~����Ӹ�ԝ�$�lyj.�TV̓�W�;gމ�jh�|��/:#e�t&f��u�.7w_rH���IM�ёRu�a\2_��|�:�Y�L0�3{�k���h8iH���]��a�A���o����$	8]-�O�w�O �|���SFmD����PL��K�U��c�W��׃ I��a:=�h����v��t�5��eȑ����g���T�R3�7���K�?��T�A��PF �z��� �6�Xt��H��v<�(gs.�9
�ב<�ڛ#܇6x��m�I�_��+!��&`A��6��D���껬��}fW#������XL�>�t�)?.uf����2T\}ϛ����u�W�[��� RQ6�C�f$xXlxV65EB    fa00    26a0�t�]��
�K�F�%���:�w�����=�|&-��Df����ef���G<���/J���t3Ite%�"��i!LE@'?���,r���a1����j�^'�]��ض�|�/�d���J�Fo6j/<*&�Z�,	[���x�l/bgX�ic?�|E����Q�:fEelm��-a�C���(�i�?!�Ϡ]�_�F�\8�R]HӍ\v��f�U�.������O���Y��.��x�1p�Um�irX��\ǉ����8Zv�����B��lY�,y&8�W]:-/(�����X.�y]�_����HCX��8ZrgÃ���{`���F��7��J5d�`Ǫ1S
�y9$N��w�q}��tFk(�9��FFq-���v���$ε
�h5�G_����=���t��]�g ��ԉ��'sP择Z������?�(z<�h�:���AZ����G�f�0���<�F!ě��#
������6LC�����T�	��
�#,^�*�Y�#��E8�r|^�u\��Wb������B����1���[���t�u��$��p�����d���;4zl/�6267|�`����B*�C/f���,�W�'45��Eǡ��y��sU����"�X,vqǿ�����7/�Ͽ�~*-�j�6XP���>귎���N��͢2���L=ٶ`�V��Ne��ڄY9�/+���A��@\ې�B�m�l/�ë�T�%Q.�`�GӍ3ӱ��N3x[>C[2���Xe�@H2v�!"�U`���|�O�% �#�g���.��~bq�	ӳiX!�����X� ��2��i�#R$��-���nӴ����ޮ�a��,���j��?&Xs�P}]�a���$�����y���ܴ?K7��U�L��'�y�:�l�Z���hG�U?�������B������!���O{���<��\�ES�=s�FA:A����4&(#��jpSx��ҽ���Z�j�9�U� d���*�S��To�ma%ѹXª�,��
!|�*�͹�|YF�@jG���|��e�6�{7Z����)����ቄB��p��7Ћ�AMd%��8.�-T�	s�=B������`��/�\���˅k)��4)�|���T����|�W�XMg�~_�/�0�0�dϣe���4�Գ1T|�4ר�_"+�4�!�@���>��dt���ؑ����v����p����S<�ǹ�9¦��LI]Ec�b��P�"�M'c/NK��Z�����\`�B��I��q�i����:������J.�@��w�.�e�(�H5��Z�<����s����C�'j���x���#�X�BWI42�U��`�w9;?�a�e� NiM�Wx`Q�0'�z�������o�����B]ic�W1(̗E��#!P�3s��},@)��xt����P�+;;�|}���z`WG ����w���ǀ�Η���+���� � u:�.N�\�`�{��L/��4�ePuP	BeKc�� ��FJ���Uq��9� ܟ��>�'�f3�_�S��M�)l5�`Ye>��A�E?��I�R,�v{�m&�ϙ	1��R�}T�_����U�>�+hٯZr�S.vL�Vz�����T܎�����2WFl��T�Pc�_�b�:�&�V�R�n��S<դ����-�����[���}��f���=6bfm�9���^�oZ��)�w���.[I�=�@")Y�5��>��;��`�CR��U@o�@1릪��]���]���45}��Ö��O^}�s��W`0#(��X�����ؐ���a�v�j#�1�
v_��Nw�lΰ��6;3�[�̀��-a@�sC�I�'��.�򴻩�v��A����b����@�tb�'�jL�䜟������S�PQ��锁����S��{d@?h����w5�\D�V/>-C�]#�ʔ*� ���fd�V1��	�gF�����A��<���v�5�H�5J�_���5Z�
��\9L]u�N�䛕�¨�*�#�� �㡎	�G��@Y��)�O��o�?�y���-�2�<��C_�y���W5G��-�����M�-ӫi�s�� �cOl7��1��׹Q�J���>"v
t�ϥ�NZ^#{�5f�;�f2��ԋ�a��J��헬�ޘ���X����L����)H���n+ c�U�h�����^-hJTG岺Xs�3�����=��;|���$��%����U�$�@�,��"u��2'�a�:n��+s���M��\+TA�Q^����[���Y�ܨ7�J��� �&�bT��s=����"@�(`��K��v���0h7����k3�V�3QOw)B�"긺�4H���̈́v@,G ����a��9��mOZ�����M9�J��,�gG(}��H;$�� ���f9�t
1S�8�ALN`\u�� �EKxg+4��p�.׌��-QXAY.rǑ�0�,�H������/��A�X�Ǘgi0�kD�ΐ&$|��&%��e��)�ۜm�痓'��H�0��t:��%�+
[55����d&���O�0��`zmG3��.�w�ӌ/�4��r/��Wڹ��J��f���@%O��8�B}YT�M���(We����#&����,��Y��F/(�W+9R9��kκ��{��g,x��mF�M�4���_���N�Rg��pG�ds�E#-�0$XN:�[.3�	��w[�e����z����p��SSt<~���o��ĳ�{��{6Ov���k�ސ_�dp��2�.�"�40��E���Ԝ~PZV�lX\B�I���՛2��%�Y�����<묮��&�Fg��4kK$s�i¹nJ���H���Db:���ǞXħ�Y�Մ-n�^ʁ5Kl�L�\{<i@�R��*�F�=���Ɖ�0�Z
[*�NW���e_�����O����OB�C��.��)�I�ȡ}��&��vlY��)�D_s��&q�G��ۘ�wԀ��n�	Uu�9��^�r�z6eN���!�v pF ��Ww3�&��$��P���[�55w���۵W�3\-@Pο_UF�d��t�$�vE���x�]A>�Әf�#hxC&����RZ/�ʿ
1���VT�7�i�y$$�F��^i6pA�TcY�ű/�#�yJ߅�V	��Sx{k��H�W��[�m�N4��S뚂'��ov���|iয��M�oUU�� hF�/�˻����1$2�b���շ<�������^����͌$!�T�ɋ(5�3���N����Vd��V!����\�2rE�[4S��NN���:Y�UtzD��v�ZDbס��p�ݮR�ⴄs����O�<���4(5?b8��0�Y1A1��u)�/B-y��s8�>F������Zn"Y)������������Z2�=�_�������?LB��g���f۸ۍ�������<�u�xf
�g�9��l�*5cO*5��!/$ava�t_�7RkFD�V�`jP��`���L@B3�2<�LMi!���qN"]�������/�C��D�/�n���WPƞ�)����akP�7�a3��T����b�*4?��h��~���aӀ��[�H�{�xƭ��:Ol���%�0��.��=+UC�6�P�.3H��[��n���f��d�O���@�ܣ�М4�]���<-GB柕7vV����"w�����#������^�G��*(�<�r�JM�X��|�$Y%�Ǭgjz�-�ӢmJ��V0���c�k&]����\�YlaYP��?�BQ��n����(�\u��MA��$�\��]�fe��j��N����b��E���m��簳�]W�+�V?�eg�<�̫������r���ir��F��ƾϖ�Yѽ����/���[�7����1���x$8A� ��B��֏p�E��T�8EZ����d���K�$S5�[�`�T�����ebc);Gkt��2t�9�I�E%�$|�q�� ½�����n�x�z)����Y�F ��@ƅ*��B:��s]j6����$�3dz�@�����˚V�謥L�zK|t����;4�f��~�n/j<k%�&�ﶴ&��?�&!��G�-�cn�s�E�����R�ܩ8��.���<vCQ�Nq6¾�,�;46g�Ĩ�����죬jR!5�gW�,����]��r��k��t.�"��y^��"��1;G�$�<����M21k�yرr��S&㸈�/�.Q��������m���~�T��['�_�X���|����cbə8�g"�ۓ����y{J~�����_����ۀ��1�~_��˼/4v��TV��9��4<D	P��L:��I�(�@��d+��S���oA��DY�_7$��qX�I�X]hqG��z�k�.�������#���B����%?�}�s�v�-��ѧ���2e|�ֻ �ǙL����I�}��|�B���)�:X	X��MvOZtݸ�+P&���l��.&l5�җ �Q���G�
�uE�(7�
|�?�$z��R1>Jˎ;�T>E��x��(Л㠵q�,�E�
8��"ǧ/^C��J��/�5��&�x��%P_��n�qu:�'�%��o��}�S ��疪�D�@�m�G�}|�������5y�*cl��6}�)��I�m��t0���E���L�d�Ffȯ��ٸ
u��c��C��x��h3�9��r�z��ycc��[k���d��4��c�n/� ����T�$�T��d���H�d���s�6FI�\fZ�B(CڷJ��O)�l�[�k����m�w��c�Ȩ��cJ���L�{�Lb�!�C�VN�z�]��u��l�v����s��8��1�d��k�v|z�Z�a�l=�G�P/�sȀT�Z��賛��z�l����y�&sD����G�T�ڒaJ��]Av� =��(�Q�HCW�u��o���xY{[��/"?7 ����2�;(��tVQ�1�pm��w�!����� P]+R�Uz�u?�~YEт�r��)#�7����\6X3)=<qC����wL�
&t�O�>�����Y>Q')Y�V�;��K��ɾi@e�B��U�����q�u��܌.����� �[]�HG�6Tܳ�4}}>�����3��fI�� ��f����7`ʮr �l�ܭ�:rV�����c�)���Ç�	�ԩ�"���2h�Ƚeֳ�;�� �����R);��<�k_!��O�p�	$UC��w�M�I�������d�P��cA�D��L�]��~'x*�H��4�� de��v"6.��&�B��:�l��	����o��R��B��y� #�2�3��Ը���xQ��E+��1�D��j�����9?ċ���ϻN��hg���Σ���7n���� �� Ŷ�>�`��K���3>�>z@sa��՞靱���RM���>�l�(�N�Wf�@�8S�L�^�2*�:�����&(�<%-��sX��t��{"Ž)<^�Q<�]���*��X�=�;����7Ţ��������:���;�F��E_������Q�4��Aoށ�G�����+��˄�k[��yM�
i^�#,^e�غ�q�_zc�p6�ߡ;+����p*�	i&���0�K2Ob�w�Q����\�q��1��u�g{#C[��r�\�I��?�R��>�R;5�U�!�J^�����D�4��?��)Q��X��j�c��K0T?����~�l���.�w��s�Z�'6��VxC=Q�I�Hd�Z����TG��e�Ra��_ނ�8����K{��1�HTe�Mu
�T<�Ȣ]��g�F��r� �xÐ5�z���~�b5�n����L>S�y6�睜MW���Har�G���� �`�� �s���%�]�T4�ZG�Å���]�U�~l�;�����X,<�|���n�F�Ǳ�E�*97g�/�8�%-��h��W�� � 7�Z��Țڠ�Á����F��)m�*k��s>� 3��p���sD8����i�g�3�n�G
d?���q�=Qo�W`�ۮC��ѭ�����9ǫ@ƶ��{�:��C����)������.CK�u#�����x�h`�0	;(q�;���=�ZnF��3�M�v���~��)Q0F3��(5�+�Բ����wn�Y�����ә�k���݌��}M��ĝ�V5��C��֙�v��� N�� C>ui5o����nǳ�������g����ncb�u���,ʵ_,s=�~v�|ؑD�M!$H#^94�Ђ&�٭������A�r3RM	��e�nRTY㧔D3��e[�}X��;G���_�����ݓ,����̮X�DX��0��NCVfCD�m�*L2[T��ɼd�M���rN���|�JA�\����tS�����`�@r�t�[>���2(����w�pҹ���Z���KK�ǧ֚k �_��������t��S'���Q��>�p��AuRb�l�Z±�^�E(���?�x薭^3��sI�6�y�L�b���WAG�'H�%=M�TI���ۨ���n'��:�B�9�#��`�:�+�*�*{�*2#����IO�9$�a��S�� ���?�`R�����@04�0�N�D��<������V�d:�Rg�lae�2�Wa�nd6Qan4�d�E��g1ƽF��S�Dw���K��5>k4�_��	u4��������a���E��(���DA�bI
�|�8$���c��]RdN��wIT��d��;�gөBjC)�,���x��	�C1�˹S�g���هR������=!��Fw��U-�)��=Ի=J%w�[�l��fPz����v�5��"c�q�VD���V�c�j���I�A�U90.73�m�U����Nb	M)(��6]�Cr�{c[��i������t�h�|��k�2Ǎ���mz�����e����o�P�3B+.��!m~:���i�՛��LY��n(E�\�>L ��":��Wwp��\��c��s��m���s6¿����+}��[ρ[�ћ<�+�R�"g����eC��l?
m�/�l�MD@;���i>���HA���G�(`u��mR�X#��c;�6*��2k�4�l4*�9�W��=�Y�.�FT�.RLN���x�K��	��Sp�eC�@9���+r���9wh�::zO8�J1���6��]{f8�K R��2͌�S���3�Q����/�����FǊ��>�G���c�5��j=�{ny������.����ߊy���Ӥ�Mv�����_ݜBwx�;�>-P�8�彘;Z�yQa�y �,ϳ�ӥdz�[]���3y,���O��j�@@���6�G�-�����
�
ס�,."�"=��#+�g����CYK���6�^!X��.�z���$|9���!�����O~�U��qE�f_N��H������{m���kOt�w�<[���t=���)�G��+df�Xx�E�s���KI�(�li���Y��
e��1�lr�^��U^�G븵���a.e0��h�!n/��Չq���ҝca��NAC[+]P��O|F�j�T����	����i��X%Ԇ2�_��iNp��fȀ|�Rv���2GwD�?����V 6+=N��l�,\��)�6�D)|��Clc�Dػz���/���0�"װD�m�x����X]E���?�ܩ�i�N��e;�'���CrFCr���@G���+'�����7�>d���
���|���j(W��;�!��#r��c����ɷoA+o�H����Fx�M+�b?؎�����q0r%�u+hA��
��tjMP�CW1��(����d���|�@�}���I��siZ�����>:��pB��2��)�L�xh��{ �)�F�t�Gý��,��=H���If��Q��t@�g����>37��nC��Zҵ���N��(k.�C/@{(����ڟ~� �$� G����8X��P'�q����klipfʔ!�2�䇿6J��k�C��`Z��:s?Cc�s��H�t�-Z��t�=GQ��$�����>tkb3<�^���|e��m�'��6�����U:���]ɍ?+Q�%��b~h�?�mJ%B�5��f���[ ED��<�w\����SGu����#�_�"Cﾞwe�z>;e:6o7շ��E�2�	J�1CǬކ;��+�q�:�a�$�o6"��Z�*����D�֙�F�n𥖣Ј����<;�!����z���m�"�]��[�*�3���()�j6��h����m��U�C1��R}@[
���=�Ј����-�b��PJjRgX�?Q�����)���*�Cc�Ϡ���a�H���E�'!�Od옎$�sC�R��q	w&2;��G z���G+D:=��NrN�x%\pk��eLLa��Ƶ�>�1����o�w;/�hK���t�ɘ�{mצ��^��2�sq!���t����H����*�'�OMA �������t��{'�����X7�)�Wf�X(�a��y�ex�`�	RE2X��m�g�$�4����C��B\":��Z�1��F20e�碛�#8l.��B���0,sH�*`�Z����L3�蘘U
��)=�%b�ӈ�6W�ܱA/���d��w��)\���l�G�D�a�^��
P7��l��L�/��p5�:��1E+Y�Ds�s���e_�ۚ?�����&dĝ.V~���d����pe�ޮwԫ{3��p4�?P�@��{�8=[ܗ��-i�"�����1��n-�X�}/��ٶE�F��g!������˜ӫ�R�����g߆�T�D��(�-�?�\�Z��%��n�i��4`���e�6HX����q�M&&di/X�����)zi�d��/��Ã_���{ɲ��"���Rtw,�oB�l�-�ܠ�Wh��v!�g�!�
����+�a��[wL����� ^Mq9�W��mnv�s4-� ���$7���f���D�u^��Y<�ZM��,�$G����\X�ؘ#<���q����83?�-����yF��y�H�Ӊ'7e� ��c�"&�&�		A�YfF/��@۴�"u�J�R->�냄O*1�P[�
�̷�Y���.����'@�2�GoތM��}$%c$�%@�����4B۳���C�^�T��7���ꭎFw�n��5&���mGI⚀��������^p��L�� 	R�G�8߈Fae�^�	>�k���{T�${p/������ƹ*^Ys���%
��qZ�;�$����@�aM;st���f�����P2�Y�Ψ,��y�T����{���!��ux9؞7EEw���<D�^'x�����r{3�=`���$�!(��}"2A��r1,]-��ykq��B+tW�tui���S�7��*��S��q�?���W��7<���E!������4�3)�m4l�~,DH_�M�;=5-�~��^c�w��Y���R��� `<��|�ix�喊d�ak�`�l�۰��M������q%�V���r%%���Έ."(��/h��#����U5����f�~q@L�z"�P��te�o=E-��Ⓜ{�S/X�)p�*�DZ�)�?�U�H��������.��Lp�|kN>�A��XJ�0�b!SR!w���g���*�EV���S�����r��79������q�x�ڿ#g`�	��yd�!�@��[3w��L� ��@�%]��ƫ(�sÜ�'\"H��g�Ҥ���1Xb�0��?J$��S����d���P)�s�t��S�4	�4�~z�^XlxV65EB    d79c    2230U���r@ޡ��@�TԬ��Y4q��)^�W�W�`^�/δ�ܞJUvf�F�ɤ	�7'�a��n>�������K�H�i6��i��&�9�;!,T���Y�[S��D��,]~-�FRL��P*@w��~�:��2!9>�k��k�+9[{9F����D���l y��'���)\Q���- �z��|0x���2֕�G���Cl�h"���cQ�r���-+�τ�HX.8*G��F��Ϩ��ӳk�ɏ�z�Y�A�%�	��+����b�����QQGiyS|@���������*��5[��_�X�/Y�Sc��W~����G��׹�B�$Q��b���Pč}S�®����E�oKBVk�3u��&�g|���>\��F=��m^�&�!
��H�h+�Q`	�F���D����w�F��-e�ZWH ���{>ȫ�=��S'��d��AE6'0�8��A����h?�HFF��^��C�xĹ��=���JA��(X��8���ߨcT�ޝ����4� �ؑ#��(�Va�^��.���{���Z���R���[.����O��IL�*3�11D:�ÈԤ�iq)�ȏ�n*-~�c�Eq��)iϤ�!��&q�^/N�=�����檫��wڐ�*�s�j�� z5�����is!�$�f��0'3��o����$���N�����<� ���օc�ޣatc`��t���'Q4z0I��b`�l�N��G뭦�G��s�Ոf�cG�-G�;aXz3���w��;����z��z�<� ���i�n+�n�(�qx�$�;�"!���Mu�!�S�~����٫l�/��د~�o7㑴Wh�-�b.��!���lS�7���--S�����eA���$,$ fXd�f	%Ut�|�
Z��\бA��Ww`2�o�?������7��׎UՎ@�K���U���"��N��юz%x.лM�	Nm%�1�� ��s��s�۽}	���N55��uT϶I�~�k�)ͷjd�s�n�4V�,�U�<�$ɛ3����(b�Z����c蚰�#,��ͣ����f���AݡqFT���ұ����ZÛ�ۘB���>#Eܥ�ف�^�����JN�c�����U*��`�o�	����a�2( W5��i���r�Ȟ��Tq���G� �i�0���SU������#e<�����(���A��ձ�͔檿O��d�� ��5�,�3�U��,]Oz�aB��K�;�gG��"�w�v���O:`�EK����>���Ж�*��A�.�N�C2�%/t��cd��k��J^Q�iG���$��ŏW<SExon�,�Ը�b��?};�>�a�(�{��q�)5��r
��a��¯Rإ<`�P ����YZ�
Ht�9��V�$���߾v���`���E좾��r��N�3= �G7�~u��ڑ$!!=b�v%8,͎c�Q�<���YQv�^�O���a�EU<�П���wfh-tU��>��F�C�۞�ھ�DT�7"0�Hǉ6Rp�F� �ah�\�e�+�L�Ԇю�k����mִ誄d���Ѥ�շj,������bNm�	@��EEv�P�M~Ӯ��"��6�
,�:�¶X]ɸڊF����?�>Z��^sE�:͛�1��f6�r
�m���| mKx�ٖZ��Z�a�+�ƌD�Z�H�m��Ψik�"�g��'mVWy綡��|��F:���j-��_+��G���6��o��=�3�,}���i�S����5i/x
V;�pȷ^�&{�kJ�����C͢�����,���K,{��`�r�ǵ1��u{$��ѧ��_[��M��i��)/Zt��΀��t5�F�c��>"���\0��_�w)����9K5�'yn?�T�6l��e�Y������o�ןs�c7�[t�ª�f�s)��,��gel�Ï#' �'x���DA>X�AK���C���Eg|������rV�5	j���O��	��x�U��A{��5��d��T�_d��_Yc�1	rlôʡ�sof�1�)m� ��C0F�?9ȸ��P\�r7[�^k���R�d�#Y�W���!���M��U�r0?�<�]A��Y=��ۙt�3�)�FN�ɡ[h4���-x���}��u���**�a�^��lv�π ��yP=�i���?�A	�i .��/)��.�6���x��c
c�թ]�o���lt�#f��(��.W ƁO����!RA:��C�+��myvQ\��^�B`�'	��ӳL�v2e�Z�X�IbT9'�}�Q��@��`��W�wrS�v�(/��hZ�w��xsܶ��_�(̄���=���)����r�]T1s���y�d6�5�~��%lc�P aP���y-�)q�'���9u��ἄP�����zp~���?D���\��p���(�����ͳiZK�;+��/��1Y:}�w)m�v%�p�P<�@@�[L
E����n:���t��:="���kG���>Fv�B`�s��p|�`��2Ծ�tS��%&,�E�����S��j�Zǻ:�7RH��z��~? 0�
��)=��e�hn�e'j3��|�ކk���qtQϏ��T>�e���$��0�3��E�XvL}��|]���SJ{fR\mkn�P`h]b��Q����̈́�����H�z�{�#V�A�5���м�ǖ�h8!���AX։.�+N#k�p�/M�&;/2�v��砎�R&�7�
Ε��ʰ^Ξ4����ԫ��~W��Y�Vu9�T���O���ZI���F�/�}��ˋ��W�k.8ke��T]@��ڪ6���i��я��z��7:Y�eP]�F5�t=�'g��GI�WJ{��X�����I-\�i:O>EG(X�=�W�}b$��Ύ���9>�C�⚻cF7�����MS�e@��6=@ѽ��93uyy_�?P#l#_�mp�=��q��o
��
T�%T�"�g�cD��\%��;��c�U��Z�z����H�0��緉��������4]O��D�G���xū
[�.�oϱ�o����I�;N�7��r�@�/_Au_�ӻI~���ɧ"���@[��Q��Uw�~�I.�Z�6����bی/f�C��8�iA��D�<���xsȳz���2�@z�+��*K�)���QC_�"�$����ЯGXn,�X�;���as�NS9���QEύ�K�(R�2`/�҈��7|x\�	�����f�#�}�r��1*�e;c�#Vu92�z�Oϫ�:F�ڥ~�<Cűͷ�DKY�ѹ��Wv�)@�4Α'PTQ|�M�P�J�*�	m��M6$��i&��ü|�ؼ�/�ըhFULb`<���=��h���[Zp� ��H� qπ!E6Z2䢵Q#xRY�����Ց@18��v����=���1XJ=D]�]�l�^���+Υ�6�!�	)~�{J��@bO���t�f�2��F�f��@�[g�d�0��%��m�_�H��@g�f�U��X=o�ҭ����X��kB@�i���l+���ҿ6{��öR����&�kl�����e�5��/����i'�(�.3���>!�Q�o��$�P����]��W��`�ٽeqggLCE.�|�r�r��y~Xr�.���?�_J�r���d0ѣ���I�*��>�kM��b�\��J���C�Xd��@��d��ae����f?��!a=.Av��y�ش�'�<����CMەG��aD���,�籑�az��+�'���-% �0E-բ�̈�Y�{Ly&E�p��abb�HE�\� �Z��8	.+ʒ����g���Z���ŗ�,<<վ44������E ���>v_C��@�R6|�\�
C�m�m@���w�s��䊵��^���rS��������#V�;�bn�4^���x*�wf��pN�9��D礰�Zc���[Ix���XJ�b�'r=�j�B��0[G'\�_�Hz�x��Ж�;Κ��o5��=,�7�/{Gۥc��i��@M4L����.�%!���j%Mt�R�g�*Ɔ�E�p^nD�
~�8ھsc��%���0�7Bμn%�����ƍ��^�F��[!�KD{-!3�Mt;��EK����~�O���.b�>��3ǜMe���J��~��Ǒe�W�����l����¹(%��'�Q�=k]"��TS���#�q��s([�J�P�O�z��n%w�Yx��?t�B������F�0�y�m�8�C�lq��Ai��_Mu�'�@TC�5��2X�CA�I�Mfx|կY����l'�͏
?u^���7��Q�s쳟5�w��������%!x�®��@��k�\�7&��6�z=�_ըG��N�
C#e�j.�:,O���ڞϨ2���VpYj)U���f8�x:��mk1�����LY%Mp53U]6^��پ>���Xh+/#�YrCa�޻)��iT��/E(�-���w����)`�]Um�p}=o�W�\_��WLQT�jW�:�by>J6);�J�6DZ����U�hr뿉ѧ67�F�F��Tߎ�;���&�Dlǳ�|yrkP�	 S��)�����ހ"U��(\ �rrI͉���M�B�����V�������ɮ�5�&c3GD!�ؒ:��XQ�u^_�9� Ё�^�!�D���}��t遯͜ű ���^O�ֆ�Ӣ��͗��7�:�	tN�-�y�:�P%I	>�k�Bt���(,d�����a�j>ﶢ����?k�P���<^�Ԇo̒-G�'�M��e������Q+/��vϾ�7��������Dv� ď�b����y�h�H��aG �zxav�P��\b�-������������#U���(�|�Zo4m�^]��Z�5�ںv��&"/�x��C=���wR�F H�1g�h�
����tNI�vݣ�������fR6/ϩhvz6w�>�`�T=��> !Ph�|IY���t-�Ѕ��ß�o�p����ui �N�?W���:���n1�ຬ^���?m�ނ�^�J��QW�Bg1u�@�Lg��C��OIaj9��N�%e�(,�v/�	��״!�mPN>���Q$���lBaE�W�?�*�%p]%��9�q����cL��&}��\YQPbS'�n^�9�����3Ps[��Q�:�<>�(�%@����껣�d���XcDV��=y*He�3QS
ug��}����ú��Ųm��	sq��}��ׇ���,;{[��$����g���LOQj�4�ݗ��8fjct��M1a�%E���5����V���OK�u��'����Ϧ�?
�"���y� @Ī� vRT����ף^?��U7��`��#�k �k������\�p�fvj
<!��\�ŀñ{D#��r$"��,�b)S���Ҵ��u��z���
���Ew�qu��0��q�����d�n��}V��/��{��u]���n�����b��4�ݩ]s9o�Qߜ�{M�6�v��2\�^��t�``���a��6�LUB��P7eF���s�o%�/ß=y���*�oEh��/��:8���W���
8r��e4k�y�اN!x�dy-�� W;��]�G}����zѶ7��G S�i��a���MF}��~ =���V����Y��L����
���AM��Q{*�jg�%���\��>�[�Śb�s^(L�T> 'A'�I���[�U-����Kv�Nz�?���%�dw�W�4��[��0���>��f=�W	I�O��J��a�ݙ:��6~�e��q�+!+S�������߅�����b��jU�φ�+}SP�h,<K�Oec�Tz����A�9�^;��w��qz��0�`_�'�l��D���v���4�m>~�6O.��RR[�z�E�+�4�J�WWj��l���S_��q�'��G�ar��~�;���cSAh1�I�w'%��r�E�9&H	mME-�F���a&���_{�%眈�2�ߛ����BX@�;�: �@L��O�?f̍$Cʶ�3ž���B��U�VJ�֓�0��5Z��g�Z��E���T��Pw�n�
48~W�O�	�gNYD�"�ٱOk��	ߒ�e �K�mI�y���^�8S��Y����]a�~Z/��P���a�D�h��;���2�^N=�o�k�IR��G�k�%�i�S<C\HXILo"�M�͋3�vn�Q�] �y;�2#x�̡õ�Y��k�	,��s;2��٤b�|H|��7�3�A+;O}��v?��K��m{6��W3�޿���.��ϱ��v?��W��̭D�\�~�jg]=v�(4#��s���NFQ����9� � 
�~T!�ۄ�̉�9�W~�9l�^��ԝ%����ߖ��C7��7�������p�3�l�����דL�8�Wȝ�����ҚSRA�B/�Z��0�k�9ƖM��.qc�}�3.\��v��,M��w
^��h�n�͸�ಛy3nuEJ,c�O-���u��p��W6��mD>����vΤ�H���y&Ɇr�gݭY�~1d&v
�E���*����&D|�a���{o���K_]�ʶR�]���� dD���>F��q�@� �W>�]�sɰ�a�ہ�����%�cX'L��Zx�z�������S�r{��Q7�	�S���i���6�r�_�RK݂�y��/�1@�ѯm�:�V絁��R��H���%K$> �t�c�?�})S��Wk/���Yg�(����Ҿ���iw�1f��EE1�"�(�;���"\�$w���O�
�������f>"-�T=��T��]�C�&�S˵.ǔW�O�v�~8�c���!��V�����%�7���fR��?���F�yN��GQ��3[}��R�qa)v_J�v"A0�2�� c�0ܣ�ḃ�06v6&�_�~�eEH���0j�1�������78Hޫ���Aշ��-
����P)�RH(Ji��+��ð\lU�_��+�>Z��|~8��vD���_Kn��z�.n.�3M�J�y�6c�p~t��9c<d"x�tP-
{y\k� S�W��7@G��Dr�X�f�l�$̶ ���e��飼Hj*2�2ߡ�Uc���Oc�0���
}[w;GH3����{-�E��ַ����r���껱����ר� �v�yc�K�5,�X+�u��IO��=P��gi��b�-'���,���|� ���sK}hX�h@KɺN��D,-D���é������+���=�a��W,)����%{����� a)����}$E�B�iu�>HXb_ۗ=��'G\W�~	��'�3��{cW��-Y�@��
�9�"�!mH%v��Wktk�dEHc>�<����<,.�k=�\��\9�;*yj)[3Ĕy��*��iJq�q���UQ
���8�ϫ6�y{{� ��N�;�JY��<��d�-)1�2�������q�Q�>k!K��&x���N���aC��D��>ၚ��@����zXPG���$ߏߺz|����y՝�!�=�L�@x3�3.���Xi�kI�;��(Ϯdϋ�r��s��yMyƋOX�R�O�O�$"�y����;��Q�m�t��y/�4jv�)lm�ߊQ����n
��J�(S�#�2��Y(��ӗl-;B����X�CH��OF�����z��Y}�*�_{'�h���(��}���~͹��O��O?��-}y���2��S���<����v?�tϻHH�46���Kg���%�&m�H��9_D	�&G���f��LG� g��z@��\�V���C`ߦ]ئ@r���/�T��S��P-	b_J45��:��֞�c,6��;÷=����3�lW�3��ucە�l�5*�E%`)�|�<S����#L��ٗC���S�x�ӎPxȣ�g�~�^�Z��-կ��ꔏ�5ٶ1��S���^Uq���Ôn<1.��k�n='sh�aUN'�- p��Kn���:�7�")ٸ.~���P+U�'%V��σ��$&��_�KQI��	�xyѮ��s�Ǒq��&�F>�6����N)�~Ɂ_��|�|=Ĳު��;�ŔS�� ����f����2�����<X������M�\q9���+Dm?�$���}��&�c�XK$�(�{��@7H˃klå�p�3���2�0����w�A��XjT%r8q���d&]_k`����b7��k��=�v���(<�x�����׏u�L�� -�Ŭ�RX�ƍ6�A%�{�.�b��1ݽ��m(���yJ�#��I]F�t���zj�[�PF}���Ǉ_w��dhTR�KF^�)>���Ȍ��ƻ�����9Y�>2p"�W���x�-.��I��$:Y�TF�6!�?�c�G�97���씘NI	DFPj��A!��J��6g�e�h�bv�8^�����E��R�_��
|�ok��J����v���X�DS-"n�L7��y��W߹X��U�.}��!;@�x��=Iy�4
�1M&��w������)@6�%m���xgg�[(�ѝ�F쫒w+�G����E��|��9T����������w�}�Z���N�K�>���q	\�_��,_m��,<^���>�N�m���حm��@�t����s��!�/뿔
XlxV65EB    fa00    2ef0R9�ֽ�7����,�BTƀ�A���KK�/TD�̉;Vy��J-O�y���� tM2�H\�����Br!	�0�0n"j�Mu�7��.�Y�Ű���� ����_.�1�+�p����=�=�P��[Ab�s���Y
��0�=I��Ȫ���=�n4r6�^K$B��e4���]�V]��탠�X����লu|f&�fs��t�v���©�y6m���rf!���'s���T��)y�,�H�֘��>���v�:Y�X��F���\`C%���"�щ-�͹eآƲ��~�M��j�o�M0�2H� �& ����v$\O%� ���ECe���0�����D�ݼ���
�u!�+fEƙz~!־>���5�K(V�bibͰl����
�()(�+!�,j�Hy�#������K߶ �#�Lu|�POAskP�Lv�dp@�c�tET,������gY�5F���������3.ҏjTAB��Zc}��X,$��P����-��I�8����9���)�Iǁ�S�Uj�� n�v�>�D�2e���kk�T��_}쥄y_������tkcd4�#�`^CF>��-�q��GC1��FwQ�VSO��j��ep:>���Krj¬b�Pe�d��Ly�ZΕ�s [�)%!�^j��1M`����b5⒮�2�h��H�Ȯ�����[����[	PW'G�8��Ѡ4���j?>��\W,��W�#Yg��WsZ��ͤ��U9�av����rO�)���&H q�B��:�8sD@Ѽ�[ܢ��˭N�C��R�UH��y^˘�
`N�COR��{�m�i;j'@���I͌�z�)%��r��'r�VVn�T��U_>ڝ3$���{�W�(W�u�]!Ig�9?q+.ff�e�����s����.�����䅜QY#2�Lxݯ�����Mke���r�7�Q�	~�N��sxS�6��ٝ�J�ɫJ�S^L�d|/���@��D\BiY�S���6pM���>�$�ۼH��[^5��^���'}7��
A:e
V܁4���
k��/"�����xO�W{�T�3�:�������Y�ٳ�ǩ,D{[��x��]"Jj�Rƛ�]l��(��;���"��hv��]X��$���)�[Lalz�K��0�*�^�0�a5*�It�������W�x��U �N?�K��|�1{8	c�L��x�?���GLF!dL^ĕ��~�k���6��Ԕ76���6�D�)�ݬUk��}�ND�6��W�Xd�H���87��y�i�]|�S	�H� ���&�Y�6��lκ\��{-5<i��օG��]r�L�zK�j�hT�>.$@�O�C$�߹ZŁ/���Mޓ"�j��[¢t�e��������du��迉턟�7VD�Xa"*"�0<~7�j�\a;3R�IS�����U�	�r`��q���	�/�g6y4QvD��$A־�+�γ�4�t����?n;���i{�p�`�{��_D��~H�����D�~��߷E���g�OV1ߵ�,�;�V������p 0�D��ͻ�"�V�|�@�=El�*L���x�R�AJ�7��2	׈��*^b��g�%L�R*}s؍��,�P�@#=`y��˃�Z�F`��̲��&����{~3���}��6KJ'���8�B3}��D-�Ni*�x��m؞�~׮D{EMr_�͐�u�U�F>�fxI��ƌ�q�m��p��0���ɨ���5�x�\�<�c��ǚ���bl�s���>x��_a�E��9}��ߙA�`	�Gkv-f'�j^�����Z�Y6�;�+%����^�~�K��>��cMOg*�����2~�5�n�K�a1�U ;%e���S+w�����㉽~%	,��"}�r�x��n	�XdL��ɋ�=P��;R/�iI|8��.){�n�� �׎�8~r�ꂰ���V�^��"YVhb�"`�,���DN��ܘ�f����[�O;s�I���=�uò�ŤM����>�V�t*��ڙي�IV�ŋ�t)�	!��=a��?�!r:��;1����we��zh�Xk�Ǳ��N0b�#+������[�ㇽB�u��O�װ Pn�m'?]�W��W� ���(J��
N�Xe��'���ں :>k���7�LCv�P������V�ÊΌ4��h然�����3ݯVa��~�t��b��ۻ�!�	����m}���p�!�Q��h�\L�.6�g�N5����F+P� 9�|v{�}.�22I��H��Ka��qf��:[������8V�����֮,.�Wްaڗ�� $W:.4����M�{�*�b��N����]Pz'��+��,>8�:����И=�������BR�2�f�k1ȋ���B֞N�3�fi6q㈮P-���[,�
Ġ�|V<��N�H{�%�L�.��^���z�+�k�f�v��+����V�y�yB�m��Y���t�����l �t��(�M/㴈'&P�{%b	� �oa�����v@:�=rgZ�S�e���ir�D0�V��f�x�>��w\SW#fYc��i��n*�<+cq7~ƸM~\�wjvNQ�=WW�����4�Q �y��H�����Λ<�r�3EY�a�����"(�<��BK��V���a_�A��2Ɓ��+4^?E6�pR���=�#�FY̰n`��gT���ЪΝn��o�W�Y�\�-;�&.�����ԅI� X�}�OY���![a{�O�'h��M=��՟4O3���$�7�XE�0�25�"H����x�W�sc&���p�/๊Pi�ٹfaR�(4�\�!�(K�3�vu�D¶��.q���]�X���8�9�7�(��Yѵ	�Ws"In�J)����d���@�7�(�ϧ�M<�ժ�YV�oM�j��n�^r�Y�>�lt�6͌ �����sK��ie�D� ���;݂��s)[�1N|З5�N@���v�lrw�
��Z�)��\�2s���Ȍn\����O�P�0Ċ���{���a�j<�R�=�Ӕ� ��X	b.R�A��Q(v|.�qFŕEZ�u�ps���-�D�}�v�Z���=��i�Ù$hp�vg{�[8�����c݃?���R�t��(t��9�PR�W����Hy�<;�Eb|S�?4��x
��������\�xo����I������}�|
7�`q�lk;�1s�é�։���'���6w[�t�|Ε]�ZC]�,��<���ԑ"0 zMR!��u��[qql�=$g8��K���p�)�"����@�H��ܿ�#�	o'�l8C�5�)�s@�H@܀zJ�Y��|E��uk�D� 5��N)���kJ[g�{R���)��;���/�����1��֧��ݩvةFќZ���O�!}���u-��Y,��y�\nnM��a����O�M��3�yi�^-�ɜ6��%��ah'�`h-%/�����F� t��i�:����bK?�o�G;�`�uKJ�ܦ2�}�&�N9���֦�%~�(@�rD��sK��=h}s��vKLF+�}[�}<����Cکtg(���۴\b���//�41G^o���'����Q>�
�v���HI�s2������m�0  =5�_�U<�Q\����������4��������O��H#�c������Y�@�@h!T�URQ�G�t�@�������Q�K�M렭�\�3��0����}x mB5(�T�߸�DHdc�8�X�x�ȓ���c��I�v��N��.@�P�iiމ���3+u�_�j�j7������+d$����mb#x�iC�b0`u���abm�	�'&�a��G���W�s� @&�Rl��y
@k�k�.\5�P�Q�4��)�C��K����K�i���!�����9�>%0j��/�NGJ��yw��l�&�b"��������A ܡq^yZ�.\91L���y���w�WƜ�O7K�������$�l�Dd��M�Ko��]W;k�9ґ�݈
@w�o��&�c��|e�ݘ⤀�����`�a4R�	(�; �*��7�?&3�4�eA�)��+cP�n�9����p��U�8l��+++u��j�hz�r�D��k��� "�����	�bL��PZ3K�
�K\Z�v�޶�'���{<��ގ�0W�i��&�3Ɔ�]�	Qxp_˺NhG>�/~�[#Kp�O�UE�V>a�;�^�C�|��q��`e��嗹������֨ �X.�
q6 ��Րk��<���b�[�r�e+tb;��D�T��ŻId��4V"�w�����Nu���0lڒ4˰�Ϛ�	�v}J��&Cp�����'̝I�_1�MŠ��E����Y\f#q�2M���ﺓ}%�=���e������ϊa�\6H��5�l�gN�a- ���\���]�rwR��Ww��<7�Bh��}���pʨv&bG���h��A�+�*�G N�2�<ZS�HF.�ɛ����q�Nr������S8i
���i��:
0g@O��O��Yz��nV��m���A�*{��2e�fzJ�&�������εd��(���%Z�ɵ�	x	�����Zk��;�Y<�BjR����i#�ݘfN����м4��������o����f&�*�?�qC���f�C���TOuk�i���UE%:�ķBB-���a����@�����`K3�HJe�-W����0w�R��92v�vPOr����V�l͍:�d�Հ�.^�;������7�d;vf�����	0�������9A�^�����?�)��$%�H�vqh�1B��is��/ᵀ�Q�x�C��.��i�s�!^������5� d������1׮?q�u�d��bu�/��խ|��r5"��I&5|�{#���2��!c���U}�ϟ],@�������V���ˠ^+��d�
�}-++q���AN!�������j{P]��sc-�Z2I�O�y�c[{�0��Q@��XG�FQVG;%��yp�
'�S��8NR��#".�؈�P������m)���*��CkMżЛ!�2�W0>��,^�=�k�+=9�:�Զ�@���L�@��ia�X~b�F_ny:�����)�IV�����3/�X9�IH�� V��l-�5�تѵ� !ٻ�N��&>��m3{@���秥�8��:ѱ�C0nδ�G�`�� eY*�ak��
_`W~�됮Ԝ䏯u,�:Ǌ�(�C[x{���~[sz��;Q���E��fO��px�i	3q�;O�q`M}&sKm�?:�� H)��]'���򦉽q��E�ؙa+��WJ����L�]o��a@ܚ�1�����|j��8݉O��0�-CWǌos��ܱ�D5�t��`�u�2���<"� �/�EEdG-tн��>�;}A�#��C�cA�4pZۂ� *��`sXc�fm"s�̃��J,TYI�|.<W:�i�4M�4Ț�b�X�0�$SFr�����*�&��
��r�O%W���l��R1�	9RR�H���I����7��p� �,�"�Q0��B���X�6j�㾹�?�o�IxV2��];����>Z�eQ��SѐR�y��Y�A|�L��n�u�ʂ#��K � u*᠏L"��Sl�#f3W�"TX�z�U�R�3J��%��^�Pg�veF����G�¹>�|ьs���c�E'0Z�#S�k}jV���]֫�)1�_�70��Ru������O/����F���u�,Mu>��oܹt�ލ�tP���{~�Ihaq���`�P���:�bl�<�kbz����q+&�]|��@��'�H#`q�����X�B��������9l����u�w��V!m�����flyM�2�p�!��5y�ȣ݌s�)+,�X��ʒ�k�y�:�a}���Y�����)��N(���04�w�d�گm��h���ۧF������)�������<��E�"#���9���p�v��5<�)8��9�O��vF[	���ba�	�����Ŭ%L��5�vh��ja��_t�dǿ	��2�s2�;c lƼ��h
]b����Cр��,�!��_���oP��k=$z��bD��2��c	i�ty0'��!n@�6;�_z���k��ҹ�����7��ĜZ��~�����-.����	��3�qh�j�N���ߢ�[�u���p/� �'�t����	}�8����_��|u+AZ��%��v�uKȒ��������K�"��pZ���}�C[���;��F-����]�o#J���x���K(tϒ�r���*�1:)'q���Ұ\�#RR���pb��[E=��㐴1���O�$��{c���R���ۗ0�~0��Z6@��s�T�ϴ8bd�2����(����$�ϑ�qd��q}���+\��\��ά���'�j�Ȥ�_�߶K��+ZxpFo��,k�'��r��b�ň̳<��{�����f'�̠P�t�p�&��6�xM����+WpH"L����O����'W��Ze��ME�o�ܓW�]�9Z�f{[��3`i�h���PYqؼ�!��~a1n����i�`m�`W~�����c}���,�㘇�N��5�r���q�^�~���/ɖ�G�/�a��>j!"^`����$j8E$�.w��2�}b5�'B@�t.�LD�����)�Qш�7[����=P��h6(R�r.4k��D��W�;��.*�3�?��($�a�\In/g�O�ݲw��u,��7�ZWWj���o�G7U��i�da<�����Nv@���Ka���1G���KӮ��i�ʁW�r����P��<e�X���I��}�.�n��m�JG�G��#��l�-�i��l�-�5I+t0̗ �d��ܔ�Ji�c5Sb�i�H�n<V
��-B1�w��5=� �������kb�23���,Z`�v�d���[N�j�V̡x�yAt�r�!�QU���5\��ܒԐT���o}�Xk˦^��4KR�GsvD걶e dwI���J]q&u�Ո&	=��ML��i��	�,�w2�B�L�q��{�E����*T�Ͽyv�_���ѣ�+����n_�ִ�T�|$���=R$��eӆ�3�1ae9��B��.�H�����_���1�
pT��}?����p�C0�����qj_YM
Vx`F�Md��c�u"�&�s�w.Y��%�sd�W�Jl�O]ʟ������t&�i(վ'��۷�����]0�x;�й��;jw�x��;V��&�Q�g��>^��[��m��ɧ�)lT9�.�$\��P��ӑʪ\!kNC	Π1�J�l���0ݨ~�����xf����'=d|����ZK啐\��/]��<K�Yz�O5��给�g��=5TA�A2�|��0��m��T*ċ�!�jo�e1�E{NE���JD��ꋭ��u:L��͒�?�6K╄V@Dv�\)��&{7��-��Y�Y�!�S����i
�uw�8�i�������/���Ta�y=c)��*����ў���5���5K&�Swb�8gS(Fw	v��gk?W�kq�s���.B�&��#�E�%AŒ{�.&zߥ)KX�Ke�`pک𭙆��>�AݓT�܇ǫ�%Hh� �v]�����aD�)�,H�AՖG]zF*�N��$xJs���&0�/��:��$o�4��Ip&�!P( ���l�H���j�뼗��0}����C�r��I�{5Q:�+D�~ﱃ����=�X7�+ycn7u�9,���#�8�1j�����q=
���� �}�e��]�r�ɲ��:�f�Z �3
��.�����3�JNB�bI�������hpĮ�՗�"8c��A�Ԑ���X���|� �*�ך.[�
���}�b&���Z��6ёI^��-5*����
�W��������>:���koݰ�����2��y���6TaM-��Je��W�)�M|�{�V���j$Zy��^Q;/��C���c�#ŕv0M�qJI�� �YlfD��� t���*iI��7���{<�s�Lq�J��)���r���юg|��էC��Ty����'2� :�d�egX������6-�_�����4�yPV���KS���j)%0�j��}����,�e��hd�/m<l٠���$�-袋�S����Bx��u+%�������kV;�-��-���t(����[�'�����EubF�!/{�q��g�)R)��n�97ђ�Ƿ
2+)�kMJ[V8�̍hqk��l�<�s�a�Rg�>b�y/ji�G��v��rٜ�r\�b��o�G�V�����/J.�I$��	�J�m�����F�<�	¬W���t��fN���d�VUN��:��B���-Lg��3�g�����-�,�q^+����'J�������FՃy�q��U����w9�<_�^f����)75�P�qd�_d�A�A]R���ܚ��F�5
)�CTS�X�n"B�PK���a���Gu�[��7��w��q�!p��ց��~h��}.��|���*��^���H�#(˶�_!�N���i�/���� 7�����̉K��:g~���#��l~�
|�)�h��<*Ń�k�U{�PY��0�Õ����Үa�g�,�8��~�l� �K��W�a��T���q�-R�H��K��V���?V|i���q�b^�&z��ytt��n�2�4���Hp�v�n/I��M�N��o�%u� Ք";�8�b�E>-���
�Ά��y��Y܄U��ĉ/��P�98	�cN��K�j�G����ߝ��+l�A�w��"%��H�cV��PS�='�>��S�X]m̴�դU��f:�z'|5��7$"U�{�J��_g/Q��g������OD����rε�^/���\U���ٚ�!W+�$�+� �_�Etr0�o�
��K���u�핲����q������e`x��t�Z�.b�^�MJ:�z
�͸�_�ձ��O͌Cau)��;�Z��&�%(|��m�*)K��5F���mFg.�Y�@Z#H���2vi,� �b���!#��Ց'>4J�(l�)��a���c���D����a���Z%�MA4r�Y�ՇP�`H��Ch�ի��#����`�5�=���]�dr{���'��כ�����#�|�
���"��>�z��8��vyQ%6�.o[��;�Ѷ)���q�5�)<z-_ bI��뒖�:5?�dq�����B��R�ߢ��"���>��<K�Tzɿm��I4��v8%��M�t-�ź���_�Ty$Op��q*;�=��\��,�;n�j�VEC�m�zsw���*��#ɕ��k�Eg'�8?%f����1���\�t-;���K���4u�0�O�-7ཝ�=Uf�0��C'}�	���B�������T�Q�4r#��,��0%
�q���%)����Rr�߅ �/���38�2�M:��\��=edJSr�����\:��&^8����ٸ��L�p��t\�8�p�����}W��V�%3P�F��!�z��=fKۯw�o�!���B��E����%����)KS�qU���k�}9�Z�a��r����f�Û�8���	��iE>�z��� #�N��������S^�[��
ĘP��^��_&�'se��	=�p�B�����_�|C�y���-v�Z�t�p}|g�#y����/�^�.Ba[��VWX$��`���ӿ����j�j��vG�&ո��v����D����F�	���q�����	�7��є�����Ī��1"�"04�GYJ,��t$���M�In	��PC��+x昇��)��"�2o���K��)��5/U�K�q���h�]��c֑W���4Y
�I3�B�&ȶ)�YDI�S@�Uɋ��,�"��R���h��z�u!������;D����O�EG�@�/&��FcE�|���Sq.���e*�b�]� �(V�"���~>:��,�� ��3�Ѯ0���H[bhҬYV�q�_̂�~���D��������e/Ȉ�+���v�7Ӑ"є22�l-�o���#��}��/^֍��4���t��1��)-�{��oól|�}XB t����j�kf83�дz'y�D��IJ�3��
�1���7&��+�yx�z\q�$D�r��+�FQ�_=g�YǑ����L�%Ϩ�[����A�/1h$��q}�=�1��k<�������N������
���z��:��(!�/���X��A`�2��l���!b=쬡�c��ʦ���(iK
wi&��X�P�`�b��k�A�T�L{"G���eZ'��A�7��,����u�ȉ�k/0oLyUet��9"��Ƀ�H��)�zM"g	�3��"�d�r4+�,8>n�>��P��9�4M���Q	n�sX��{v����Fe�nw2A{���}p�Y�I��/a"������\g������`o�M'Lb� ������y��a
��'{j�������?j>C�f�M��b���e�7��m>m�{W������K+�g��\=,k�V{�ۻ����P] C@��@�</ܲ�7w:8�pg��Ӣa!F�o֭�	�1Mk����ѭ�b�j��.˾��^Z��,��g,��C9va����9
��X�;��f� �OO�yÁ��~�8"���2鲧���H����\��'�u�B��y0h~F��X��%k&���� ph=��g�g�e86v5����n���>Y	��j%�L���r�,�o�"�vɸzY�$�ɖ�5��PM~�!���e���H��+�*�v����b\]��H�%2�ى��̄6u�i0�Iͳ��y5�5~xd'�1�A�n�c��R)�q^�2.t?P��� �3ǘ��\�ui��e�”��߷J�w!e@ kA*�ƛ����ՍK��6d%��� yf��
�̽�S����f�4� 6�"q�����A��!�N�����@���b�B3_��աA�!ؓS�:cK��6s��1zi�pC#�%|����b�ߪu�ͱ�����a�ﲆtz;��O]�=�D�[_� �:��|T�#g{" ������ݬ��^8G�N/�Ϣ-}�����0��8І�ENPk���D�(���^�>�G�py����X��F#1��qQ���|m/a��m�����k�QK�ܫ�$�	�:��Iљ���s�ڌ^�/L@�^�d��)Y�����v���"� ������Г��4,�IsD��v�Qo��,)�,NC�,�r��
���^'\��#��g�W������b�XIk���]��CF"y��UOsȆ��$"r47�ܵ�#�w6�b|����[NԫG$vclo^M�[��D����6���f���3�0�<@���+OY�SY�Wv��\�b&`���'+��p<i�����z��JV]���d���f�7x�R+��'}�$-��6�*D�B�P�+�>��&ؖL�ha��ĿF�>y��4dȠ�^3g�P�{����od��=��{����uE{I���)�`&^'b�=Y�@��I�~��R�2��O	s�0��)��%Tz��+�bs��qh�g�Z"�}ҖP3 ��k-���W�=3��a�		u`.�e�/g��VV�� BّSP��ҟ�S|��G._@��h��1���u�b��0�M��d�[0�j�y u����h��1C����ؘَ�� ����a8cCW�-��Aɪ��OZj+�D��y78h3y�"�l��a����;h�J�´C��\Q�g��u�e�l�]c�;W��k��XlxV65EB    9737    1a20-��;P[������xy�ޥފ,Q��[ꆀwk:��T'K���ft���'�@hU�)r,!p@�$4#-����I�-G]��5m͵��ʹT"��{^�j��'ړ�B0�北�X����h����)u�Y��֍�sp��f�����VN,�(�/��W�/�G"�'�3�Pܠ8�h�'����`;�6����E�%d�yį��]-�Ax
j�I��R1����������E��um"���W`���AHp�EI3g+��G����=�	q�i.ش�$�S�ogߺ׌D�RV�p����A�$���+���԰0������L�����({�?����g�Ds_B�uV�{�`.q�;����&��h�����Z'`���ӹ���	������<8R�}��m 1�z�6R��b\5�̍>�T��CHY�4��!�X+2JU�k���E.��UiP�k���6]!id�.(S���x ��=�>*��2L]�� �O�I{HeIR˪K��RH���ǝpo?�9:Xԑ�1_����S�Un�`���qVa�����#� �ي�ݑ��W�R�Q^Z<���������M�r��;-$�qM]E:#WL#����W�km �tb}�n,�b�#�f=yt�n4k���O� ��׵<�di�l�Cm+9K�V�	5ި�j��F\h������F����Kt������2�:N�H5�� ��;عC&�+�\����x�f͢�m�����-_���.O����Q[����]�\�ی\龔D.�+�J�o8�\nt�����`9�����5\��4���
�V�&��
Τ�6�����鼃f�0-�|[�jj�������ċB��6���g[�2�C����y��9u��bޮ�D�gϚ`���f�nC�ﳄ�<�`���B*x����r�d�������E��W#��ģ1��A�f߭7PN�Q4�\u�GQ��]6���$UҒM>�b'��W�S+B\����r�𡚑�(#h#W�j�k��lx��g�Κ����a���ʎʰw��	��B��g_���ҋ�}W���^�<c$�_P0�g�X���vh3�%1�l�y�`�Y�)��:^mN� ���H&`Y'aB�y͙�^F?_M�
:%o}* @�s�_؂$(f��[8�q�쓽Ɓ���?帎�����c|�D][LTd��pFVi�{��*B��/#���'���5�>C�\�r��݅�'�M��v7��_[�G�XϮ�s��[_����k�1϶.�t�����x'�~Be���1��Q��X @U��ifx��N��V�V݈8(]yecK���|�A b�t����C��U�!�aǨ}�rk���P+�7V)�����{��I��G�b��&��6���U��KH����\/	�a��p�}	�F�ȘZ�=���IϦ�����¾��1����>�Ի�H]�~K�Q��n�*p+��:�	~��]+r�(��ړ�4�ag�_k�:qF��} A������s�B��A��GsN���������
�`K��ro�%��7t�	~"�u��x1#�&z�?�l:C�"X��,E�ί4��9�����(��7�����2�	7bKoi���P��N�z�#
����j�/ ��&UKh(��5q�8��ԛ���Y/.=S'Y%����y]�p�"`���s�bљ���l�N~�|/|�_�|����I�4�#Z;�+T�_�'g
l���e,^Z�/ �ݻ��l���ݥ��w7�O��oE����Ѩ���,_m���F�s��N��V�����B�0O~RFV�<�x��1��>7+��x�Pc2(Jy��]\��A쯗��F�#�W�*+"5�ܧd���7����+p]=��r����r#d��}��ވ����x��d,U{U��^v0g^�=�1��壦zlv󛹬�M�
���+���ڱ��~�W�	%K�|Պ��ӛ��d�������p,`��4z��L&�cfٶt+2DiW�>6\߯%���~E�^ví�6��g.�K����LU8�
E�#�k�\�^�c�C����o(,30��`�nS���,�!a5��h���v�4�HRÛ�� ��/������n\����7!Ӑ@(������ɾLD-��V�h�E�[Z�v&���U�OU�b��'��q�v�2l챺l����@�"�z�z^�|�T|��rq;oL )J6�#�®҈?X�݊�{�^��C��CǄ���h���������L�����񹸨gTK9��k&�n��xh<\]��=qѤ܍XG`c2��u�|#`�#�!HBY��`Y����vXr�bqk���֬�ɬ�T����E�� ��1����d��M^�w�g� Q�s�u�z:k*=�}>p Z�K�X3
�b~;��y�2�p:�=��w�w��i3K,���Y{�ġ�//un�Tdr�fS�&1w��G0B�_�!����|�� �&^�j!�?#7�@"Z}b���ww0��.H����V���߲�:�
mP�h}p�DfbY�u	c�A�{_P�1�{��ADZ���c{b�Wh�uK�?0k+nh�W1�%�W�"���+}�����n�&(Y�_	!0KD�ٖe���Pmˉ�aQ���K�T����ҿ���/U��T��ߑ�8�����=��P�چ-���7�S�(�#�X�e�Q�ɿ=휠���@��YG�3e�Ž����]'�,̜� c�{�r��������o�
>2N`�mF+�?(���p^T�r�i�U���y��ces�j�Z�Yd��;q�������C^��3�Z#Č�{u�� 6�s_j=*i�em��M�\�Y4_��ԩ��%��p��QBZ$'�B]��fi���ّ��>���"�,��9�qt�X��x�򹞥:��^�}֘�Viͼ�w!eg��v�URL?/"����Ewيk�:74gCe�a�俈 ���+a��h~���9@Ȩ$g��[�l�K0��l`�ȕ2�*�V��Z�9�um�!���e�K��Nѱxfz�d�hv^c_^��&׏��^YI@�г@�A������V2O'�Ezn[8��'���d�*2U�9�����H�,6���n���J/�"
z�Sb��t0	�ؗOշՙ��~�HΨ*	Yc�0v�c�1���mQ�[=���剜�Ho	�.���1ȡЪ��/;�"g��a�ӯ���T���嬼��(���%��i�����M��k{�[���X��:β阍ߙ/�be�o�-�;��)�^L	ӟ���"�,��^���$ '6gm��n.�wj��1o�. �� ��,H{5����2�Q}Z�RG��:��<4PTʱ0d���G��^ll��nPH)��������M�wﾋ�����u���e((��QH^�녇��ǱO�����Ӌ��%(���`�mv�����`�V�Ɣ�:LGuD`�GW�t���п�V3'#�}��s	���_!���PfJ�$s���o�ZN�R�ݓ�v�8`_���19�N�PH�X�|�x�,�O��]��D��QAQ3j}����!�bq�9*G�����&㌧릏���\����͜��d��?J�^����I.~1�Gu��S��V[.��)���1R��l���Z���8"�
p[F���H�2QM׭��xa7#_����x�}a�":�V?���� �֋]�(�w���_^]:����OW����<�U�v���|�D��1(��؂�˙G׏/:>�p#6�֣�1�ή����rn��Y��/���;c<�t�Sy�� k�K�~e��(��O4�`� v�����qN�ʐ&��`>�t#.,f@
�L�kx�|	_as��k+6�^�$�uR�����©�� 3 �B"օҾ+^mM9���r�!	eO|㔸(��9_:$F���搡���,9�'�XL�S`Pg�c��go��������3/� 	mгfFo8�<��X�z�]�?��h�P��ߴ���]�Nj�d
������ɏ���Pm���H�k�@L��"��Uk�y(<����:Cq��/7��C/<�u�x%�KX�%r5� BZ<|#������#�*ć7�u͖�K�LxE��
�_|�;� )"$�w'�%#0�"��9�쨧�ȳ���� _�_��>�4��]S��n ���;ŝ5��ب����f��:�:�}�ր��i��S��y ��ҙ��]&���xt������X9�v���~��7����N{�ӵq�K�S,b�鸟5�7#�# 9�4�'M���-L)5_�pԯ�u���}'t1�/�￱��k����7C�\��"'��Sf��Ou��y����km��QY�Bz���>\��gG�}ʠ�������>��(�H$���~͡7�"oҁ���T��h^T��-�pR����G-]�o�@��L�P��,��&�h�Q���r�����Fq:^��
P�A�>]��5k+o�7̟^!)κ�Uj��6��C��������a�������bZYo�Ţ�xU�øZ;ѥr���jUԪ�(~Kb�J����R��,a��䁴�DRAd�z�U �ԗEp��Ѝ��0�!�oh�zI�y��BD5��6���h�F`�s��n!�F{t��	���+d����A�6!�|`�|IR�R��KU��p�Ճڱ��,�^��ٕ�>Os��:)�_�l<]ʫc�������ɠ�<�j�xۮ|�U�]��122���G��!��]~�舟����S���sM��،�X�7eK 
��k��c���бxl��C�[u�
וe�����{Z,�TQ}�\�g�����{@��|K�~�H�!B��51y�1�+#�e\�%p��*��\��W��`���,(ܞx6���]U�-7��_�wɖf�2���g�1y,��NPIѴ��J�*;������RЈ�~f�Ě}��;.��R�*�ǚ��1��a�d�4��爫�]~�r�2��f��b��,]�g����H~� �����/{�˸�zj���-|�'�xk5�K�v~F�u��P:R��\7�q��-#|پ=�i�ch��b��
���2�a9$�X�ܺ��t�`9[��v�Ɇ�@����J����H���H���I9M�2���d;���� =�*��ʣ��GV[F4�;�5$uór���t�/T�߼�~�-�������P/@ˢ��x��(\��Fnoޤ'-�F$=�bG� /����k*,�o.�3��� ���'SVڱ�ʝ���yn�����x�2Z�ܠ0J���P��q͖�&"�6jln#Ħ^���6��(�;RwUʠ���@�Ǧ:]�K;4�+��.�'�C��?wD��n���M�c��Ъq�^�@lg7��ڟM,7��	��E��e�^�]�b`K!��O9�ӟj.0��C3_����*���B�%�/o-d��G��˹�8����Ǝ����c~Az	�e���Pc���p�ՙW�Ƣ�
���|'L��*W�}E��q��7��;�ّ��|�TC�����r�dkP���Ek��#/?�8��(���m	�啘=�P�������VsD z:���Ӻ,e�(�>� �\�:<�,P>��q6/V3n�_n~9����vH�-�Hs��
���2QVn�I�$U�˗s�U.Sn0&�4�(��h�&�.���<�( 7��.����F��J|���[�K&�-���tLk��2ˑ�L�ۖ4��4pK�����w�4��z���X���f*,����8 =P:s}�������E~:M ����J��3.��~��͢p�/�L�~��En���r5^Uľ�)jɳo�Wf�w��҄�t��0�U~}A��S�/���<w�f����jbj�b���ƴÒ�%�J�����ז"?U �>8��k: juɺ4��9.E����1������A`7��P��)u���������M��Ƽ���ݐw�j�yi�[-��8�
_(�Z3��%������N)�ٖ����a^ʍd��;��`N�y�5�.»5�L�0�N�g��˶F�5q�^��˃'̼�_�`ЇϬ\wfN��#�o��Yo�dD�����JH.q7cT��b��[#��B�p,*?�-� ��j��7�ts�����zg���*�/���uVG�V�8�K�K��h1�+7	f�>��"(=�"�q�C?���[ �cU���1.���t�J ��7����R��'�e�m�s�Rb7"� �L��u�/���6H�+l�J� �OɃSUi'�c��X{�\���2���w��[i���]3Ӄ�Lf)r�^E�ee�}���Ԛ�]G�S�/��ޠQ� ls�t���mS��F��6��;q���!�N��(�V�B@jgLJG�=�}�C�3:��2�bK=|�u�l����0baC7ХR�#�+�^|n}%^@<�� ��[�to�l��dNOm<b!%�å�;�!�Ub ��; -�3�-w~���ץ���Mv�����[���OT�k���ShOH�rUL�._uj>J�e?R�s:��2��%��G��qd
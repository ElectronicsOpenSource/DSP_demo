XlxV65EB    40f3     f60�d�!d�2�����U&)=�\�VBz�_��\��Ur^��SlH�hڵ�Yp��:��gu���%`Cv>@�_�p���F�R�j�߭/����I��.�Ҵ�rA�q%�I&��iX\�R\���ɓ��
x����"��I���;�����o���A��U<aaa��C	EՅ���F���:�!���1x ?Q�i�� H0��g�w��G◜0�ύ�1�ftc��_t~!����M}�o���qc��n�ِ01,�7pҶ�ݧ�w(�e8���u����M-�F�!�|�:ƚ�^$�nEh/�&�?]��AL��1�|�=�ߣc��"�ĝY
b��Pto������W;�R�O5Ļ	Ǔ�hRyJ"!h0����|<[�Ѩ�K]����7���A��2��9.��"X�]��$'��֙�u;��$�ɫ_�*?	���^<�1�WM�����~ >ِ����ٝ�7�8F$�~��,U��y�ʡ���Y�U�gn�I�a�R��ɥd߬v=<���9�D�]IueE����'�r������w���EC���&� "g�\�����c�̐ܮ�#�d?�aj�y��#J�&��5��@���p�#��}�n�c��>5�
0���e�?JT��C����[��$��u�x]|J�7P����PF�����0&\b��c
��J�E�iO���ȇ�p�Hq�E��Aʯ�s�ݱp(���&��gCv7����9�Ʃ�$\Bv'�� F�v)��py��,�}k7�H���3T�Y�3c�o:h ���D�H�\1a�u˧؉��f���Z?��w;�30uI��ox�T1��,��j���K�8�/+QZ�l2�ч�gN�>l��f�#,�8-h
j7� ��a�&G7r�yt��P���������8��OA]
 c��.+�J���J���ņ��PH|�B�:��S���L:�Q+`�/��[M	A��9) �����^���t�9�h��� ٨��2扛|d]�-�=z�,8܂c�L-4�Ț�)�]xރ�]sz3�#��k�	��$�R������5��A����	J��RLj󏼒x��Sʧ/+��A����tI�����3$$8L����_dN�O��|��.}�.dƑ���G������5��uB �(�j���T�;��_��Lik��~JCg�=%*��q2`��e.�ـY�D�ɷ�"n#	�2�4�j�[�=�!�\=!��6��g�V̉�Ɨf)�?��J���7��mf�s$-��׾z��yha����Gj5�S�êW
��LE� E�E�dW��{�n�`S��%ͦ�A�n"i��
��q�JoOuÚ�4ߣ�z����s��&|�Z��s�-���D��$��G�]�f
Xs���S�Zj�c"����'2�����]i2�U�ѸeOr�pZ�Ed�;�3�5���'N�MP?��SV�J}(�5B'�n\�m'��[��|�uiEk����D!��6�����=��6hJGސW-��ֆ#|�4����뱑V�QP���U����y�=�Ez�5;�~�4���G]_�h���*�T��[���i��E���Ѭ6	��r��ygs�ӊ�\��٢��7��<�r�$��E�jd(f�E�ӗ�]�'zݾ���r�Jx�3��x�M��4߻�X�"5��\	ʳ��-�{���P9zySx�w׈O��%�i�[K��Y�ZS"d��͔m��,姒kH4r�^8���N�m�+��Ո��̵f�3/��r�i�Q 
����$�U��$P'�L�X*�U��Y���~�2���pU�����/5U����c�6�=N"{��l⟙�*D��s��c�r�xg���V��MR�E�����(
���� �fB�]iJ^�m�w˃ﭲ�8R<���Z5(�*H&`JfVQ�0Ρ��w-�:q���o�BE�;v�85�VNT��n���J��R)};���Rd��w���O��@k*�"SNj�y��҇�pĲ<��1���^=�a��:>�S
�RrB)���.����/����ѲdgJ����-��q'��O���A���?Y���Du�Ȍ�<N�����.�3�~�O#V�%�N+��a�N��e���s��L̢��qḱ��C�K9z����cu=���r��;*�ߨ��R�&#Q�sW*�Ƕ5���U�[LO)����(�� ��9hk#]}�>�)_�H�|0� lcgb��yԄ�R�#�(Cv���p�Ƒ!���J�V� �J��%����s���Sj���<��sn�ռ�#r���on���=��4�t>�B��Hnz�b��_cA����g��d_��uPa0��2�,bōA�mndm���,'�N���<DK����� hv�wJG�N�rRYRUtdK�w�����O�Ϣ^:���-��ux���o�E�<�|W{���EwN��QK��Ҥ2� .��0Kħ��I_�W!;pL_�~q�1�FҠ}���r��Q�t!:�Ǐ7�����%�͵��s���{�k�vO�m��Vc �b���)!$�x��&���J�K8�����v�C�ݪ�̑��@3�����@�N�0���{�L+������Z�O��X�s��<	�������b#�U4�ԧzRK"D>~}��b����+�ʢ 7�(Q!��u�j �g��G��k�z�i�Z̻��3|�t�����?\���B��ǚi���p�I��Dc�5�B/e��(��ِx�9�l�����?X�\q�u���D'D]&���T	P���dX�0��#q����wF��C�ۂ
uW3�!��ow��7�j�(�+Ǿw��g�_.(+�wi��T��} U|߁���0�"�?���p�]�R����FY��f�$���c�k�^���d�(̈́�'A�(� �(�� s�\���&H�|��AB�f���������]�B���Vo�A&sH��'��ʝ�
��2U�ˬ/=��B�����C�����=������\��e��gu�G�cɚ*`��d*4I�k$[�������b9[��Q�7���`�2��ҭ�F�T�}p�� (�(����suV	��\�����
�۵r����%��PԸ��b�r�Vư��Ǟ�{�'UB��1��H:G[���T�f"�u���q�C�]Y��#u�����Q#���k�i�ϫ��0}ȸ� ~L�R���� e<��.������}ђF���7R�}��J�u��
7����}|�B�c���}
���a�E�����pG��}��r' �.E�l�$0���Ҵ�ɠ#HM�$#�õ��o_�t2����B�i�4�0��s���~��\+�FG�S ��ര�������ʓ�72B�|=z�˫b���St�lS�k.���t�(�,�3�R�I>��E�)�#���j�*p�s�CfƫG�16��B�o�T������FO��H�+�n8Eל�m��HI�1�JQֈ����h#P�Ixzѩ�!F�k ��%:N!-)וCW�F5�$��p��:��1/@p쪑��L�滉٢�:��4r���t����7���]���;C��mXzA/�(HZ�R.����������T��޾�Vv�n��Xl�[�����g�[fV�rM�m�Jg����O�J"!�#ˉ��$��x�kJ�pZ
O�eX��8����	�:�~�N<I�J#���A��J��]�@i%pKy����J�K��m�V��/�H3�GNL�gI	��G���4��		����#��1��[W������?X�T@�m-�2ݾV��bq�XQ��} $�t��%��%��1c�B���e�Lv�D��#�V��Sݴ(/�r����t|����?=����<�Q�KU��A����#�����*��۰#'f��
XlxV65EB    19d0     9b0��!��R��=��*)G�]��P����U���<��({3�?[��%!,�d��7ظB}ǐS^��y��m��~�n/����&�Vk�HvxW���A��J&���|GG���(�s��D��P:d�6y��Z}��g�c4z�9M�������W�J��6*n"�c5�BE�	Ɛ&�G�j&4��N9��#��ƉyB�����{H�����l��@�;z\�.�����/��ߥ�&]���-����E��fU}[cj���u�_c�p���|u�Z���e�[V�W�����n���u���"y�����G����WHb��B�3�$v ���M^��##�fH2�.�7P��{k	�������ID��%F�'��JVR��
�!�:����ٻ-L��0�.��_lCdUNy8(�� ������-T�6�h0,הXC�9@0�*��V4�U�o��K�'0G%�x��XeʏT'��~狈����� E���Y����&�pц��ò�A���߯��>�H����q�G�O班���Z��ɴ�y���£P�l"�ɛ�A������R�ի;�d�& ���^x�pd"h�c�B
Y���+1��B��&�iU3M�_<�/%�pϔB n������q�`ʾΠG��xFm7c,��j�-�>y�\�3t90��S_&���ÄR��!��Ң���B�qa� �I��:�M�#R���w�d��)N�@&��F���N~J��pd@Ҍ�رze�	��%�|��"2v�29��p�<��4T͠��l�*��ܟ��&4���Z��ɆX�3T�� ,�#A�c��qa��t3��ީOY���f���\�T�����/R*�B����oj#��$J�?�}���ǎ�f|	IG�D�]J�6�p8-���M�m rz�����X�4��`�@�&;�*��;�e�p�{�%	�]���"�Z�=w����*���'�B����9b6���t$P
!�4�1ޑN^�R1�%[����P���^�1�`ˢ(����@Ł�K��z �T�����n�?���ш�2�����pXZ������/�`kl<��5�ª^�3�(RjˣORS�*�l�_��{6h89�W&��m��� e�=I/�4�:,?z�נ7<98���kΏ�h9�v�jHA|�TPҋ�0���cs�QA���7�rL˾�\��J����������h`�.�/����5
kTW����~�0&
v�s�O�H�<� t	|��3������?��������{�!� %���#�t3}�O!"��搠�T|@��C�g�"(;SDX�"L���s�m6>)�'��7�&*+���pr21P?Ov���N��Ax�x��|����[��-$��[P�}���y
��V}}u������K��B��t=@��W� E��&�Kt�(���NH�_��p&�s�u ��x�R�7���4�t�G	��!��:�\�˶��!:�NwQ ����ZD��9���{J'�!O8kʚ�
&���'��w�Oȍ�d��><��G���N�L��4��
K+�ri�I̫�1-�U�F[<\"/ݰ �U@��&.�
UXqK�g��,x���REt)]����	C?n@�+��R���n���Ӫ,��p��v��f�s��S�n����\�Q 7�u���c�?���#ے��0�\xtR�dz�C�Ly:��l�V�֤��A �_);����S)"�G/��s:ro�_t3^k#5�qE�:�t
�p�]𺊝"�(@ȓ�Gf��3+����6\`�
��hҽ[A��5�uH�-r�"�^c�|�������^� �1��O�^�}T[�5
e6칀���4���	Lg�G�.m�B��%V-���;ѤbS����#��D���d犥&�����`hn�Ƭ�1{s�kafY�\��	�$`��ϳj��d�!�m(��H\��> �u6>yśY���|���(���LU1���ia#�OWG ����kRyr��:��Ӄ$V��n�;H�B$��`��QMtА��f����3�FY[U]`}H���g��ĮX�r�l����V�}�I��y�Ed|�v���1�t��p�׮�le3�3t�Y����6�͙dX��:ͧ'���^hV�V��aCwsg��V�#��Ђ�Rc����g~q�Hu/Izl�^��K��
#���Hm��OKOe������ӥ��b�o�׍�T�X
u�>�-��I���G�ڕ��^�n@3PZ?��1��yQ`�zL�Y2�2�k��V�K�&��Z;�p&�ꩊ�=Z�~T�fW}��ȓMp�@�N�O�-�a�� c���]t5/B��>U�p,Qo�5�����r��>`<��e�G���QCCVh�.Y�Ci�,�%��ב�-mGI9��aw�>1�`���pc�0|}�`4��������n��L����4�
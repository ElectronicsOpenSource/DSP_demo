XlxV65EB    6623    1520y�����^�"�wvx_J�)�g�I@'���F"e�K����K�-�����}�{�x�/?gt�Mp0���Տ�	��(Rg������9��9��/�.,�@0e����K�����ڵ3	�]��[B�}��۰�����oO��ڨ����av	T� 7q���l���/�R�Y�&��2����<��}����Lܸ��GPp�IB�#��{�v@K݋�D��P�Mȡ���qW	//ud"�ɷ~T� ���U�v@�"��R�������TXw"���gK�]�l�1�x���^������e��,I�GۉW�|�T�:�3I��.q)����l zqP��gSzfGy|�퀩�|�@҇�.G?vв{���s��	�C*Mb�s$t��>�������a�U�SZ=~���	��Jz)ǯ�eN��sh=���<��s��.ـ��������o�:��>�\�O@�$u������VQ����e�=�;b�x��v�X��:�\��/�,�Q�$6��RE�Ѳ��G?9rz��{��9g�Q3mhT���~�[�u-?f��< ���,��V�Nf�
n�yڀ�C�n#�?��J�nv�+���E�)��O��������W�|@e�ͺ˧���۷UC�)l�P��2���V�S�v��7��d���^�d���_?���I�O�7.�ByH�u&*!���|�-]T���'�b�Џ[|�L�?�~=LԢ�a򥗊<x,1����.W�=�z��s�IVy\v/�
��b_����g2}(�|�Q\�)��\n��6<�M.d2��A�L�)�ט<Ǝ�Ӻc��6����$j3�n<2U.L2>y}g�Lʕ�m@�͔��Wr�kJW�"��4��0�v��6�#�BS����čBTЉn�U"ҵ*o$�d�ݧc����;r�%�㜭���S!	cF�k�V�����F�y}��M�c��O���{���<=�H��$Ҡ�؇�o
�Z{Ɋh\-�4N�[>�⊽^��ͭ��	��I�w-�8��,0��$�4п��g������R>~���G��Hn&	�*K��p����_36�!��ӧ2��6��l����W�Pb8gaJ�B�\s0��c����NXw�5E�ۖ �G�
���DY�Hnz9�ǆp�)��z3ժ��%���)��b�[���0��"�������lh��>.����U=g
{�I9�GPbl� V
��nj������!�Z�~�/�*�rKu>tR�T�M�K���e08��*�{	ݤ3X�;+��U
gk��4S��#4~b�;h�HW}U��]^ák,v�\(#G���M�`�,8ҕ���^%N�
+�h���=a�Ȋ��+=?��Y��T�gy��O�^Y#��$XxI�Y%!���t�R@�P�� �$8�Q�����j�<��l%U�Z�SVO��J����x�k�d�u�#�_���y��bXi�3�mm@��Ů��֩�砃���U0�Hd�����H��c,�@��Š�&,4��p�b{��P.1\Ksc������Q�.(��jC�XD ��S�c )�`hڹ-cX"}H�"��G��Tu[O]��J٠Y�G�׋�hߤr"���-��u@.;Z����/�zer����PX��H�qB������'�ƿP7���C_�sa���W�t��>W�Y�8���Y��?32�*uк���{���a���'�:��L-fy��@�������I>IVＬB�k-{\Qc�y��t�yz�b���f���gm}*��"o$�N.��{:��1�Z��q��.+眐 O��4$.xRQ�cr�V�,��>]��'e�q�\�U-��^Ԩ�9�q�3J\��2�q�|��Q�ď��Yen��:��!A����;��YYoU'gQ�x�F ʧ�3D ��I� ��Ӆ����F����w�T�xx3��E�+"�0�A�z�x��v~�NB
��IDH�p+QC��{�3����?f��:��^ ����阇pJk\2,���u���W�GcZR�͓:ƴ���Gq%�y�$9��BEN#�@!��6�8��rn�ek���9d*_*��1�����[|����e%�%)=n��#o�a���\���t�Q��O5շ����Qu��$�Y���*Η�x�R��[r��L�{�6�}���N@�Q������mi�<�ͥp���Mzr���ԑ���ͩU}��aY,f�@�2����c&A�7O���}���܌�;��IJIX����=T}}�T�;^8J�`���%�1-R�|��>(�����h	a�5��b�������3k Q�E"��~�"ۍ���������7نd�c�?�����D�T��f��{jڒ_�I��e:�{��/�a�,ѥ �9,v��j��'@�-5xaP.<��O؋畲"u)�ޥ�äCf��#�?h��gw�] ݬH"P�p�uw�iEWb�5���ϠC���,!�ȟ|�B����1MUcw��]$y�2�a� @ &K���aC�I���*;�Y�F����:���"w6 �8�87�xH�Ɵ)AYk�ȗ��|r�1��hO4+�j�)&�"�(���\�+aQ��>�G9��ҭYD~�o&��6 ,[{ϓ��\���������T��fx����z����Ն�?o�V�[TiQ���WG�$�ޯ,��[�> ��w�AI��T5 R�*�D�U+�a++������]�P �������
~h�,V�Z��|� ��ـ�J~�h0���	]�IWpEC��fK����*{"GZ��X|ě����O����}^V[7C�U'	����'����,#�I�#�����J*�!ė��t��!�y5_�1�t!%%|O7޾T�ۣ� �M $FPv�!���o��a�#��� ^r�����O�/��v.����s��֘�&��p���S(D�*C4�e�)v��P!>��
�bZ�\�j��
$*(l��?�������3�e�T� ��(*q�C�K��~�.[#�+�'�j��o<N�=��CLR/�G��D��PL�=��@
�!��#�OC�L͘{�}����/��]9��c��	M�׎�ģ�?��E���q�!?�Aʉ!�ݛ�|\�_�hŇH�X���%0�LQ������_\���;}e���������E@�f>��g���:h[j/ϻ�Ҵu�D���6pQ ��"b�ĩ��J�`\yյ�k�P�v��D�{���;K�l�B�N��p��V]w�k� ���T��K3j�0ݷ~ZCĲ,`��=Bw	�@�>v��~ⱑ�(�L1��ΌL��{�8�_m֫�e�8w����V�����q&�����R�	�4����Wx�����n�Xh8���ѭ>�R_q�'P���	Vz~^m8��T�J��kwsC��e|�ń��_&],�^]� {��WG�6�ڟ�gbS�������9w�����JY')z7��2��Q��
^�yOv�eg非}+��2Dxt�ܜ���!Ol&�����z�A?��f�J��� �b�_{4Ę#��'��˪cє�J��~���x�t*��nY�cۊ�*\Mu��HW����d��p���n�ެYz;,m�"�����ٕ2�ɀ�B"��:?�
�q�oyb�d/
�aU���ӆG+���,	��S������M����ׯ�#F�������(9�'��iF?�IC�[q=�g�À�n�#,n�˘��v��D�:�~�=������8N�9R����h������yk��s;$h��xLF�N!\I�'F��e�)sXa�?N��U$ʚ�&�}q�0���9�,���ޞƍw	0����9�~������"MX��(44��raI�
�2"������j����g�v�׾k� g�Zg��O�bY��/+����P��%u��-�6�Nu��C~�E�!�l�^��Z�#�ҹ��2������I���F��p
	��\0�ĺ$��STsh�ݕ�Ì�պ{�g�T
d�����w��z�`6Km����C�z��Q� )�ƞ�s�E�y�f�z�i����0�ȸ��~���|��v�)��r{�UgZG�:�2)�!ס�2�� WJ���o��Q4^'��М�S=�NG}N�o�q"�OQ����t��Z^�gS��r�{���Q��:��X%�O⮞�E~P�)��J�q��m�x�|5�����G�ǩm���r��f�y86�U�)�����L�2��P�`v�<��R`�3|l׀R���{�\����f�M�z��]�d�c�+���O�rL�7�� 'SF��#�p9\@�q��?�j~�=)�7��^9���UlĿ��+����ӚUv�wg���y*C��5){_qb��TG$j"���t�˫��jfb�O�=�Y�1��G�ɇ�)F�5�
��O�T{Al�}��}����k�ZSF�xt��Ȋ���g�Z����Sv`��I�R	En��q4�@C:k"V{ �zO�2f.ꉮn��NHh���b�b�火���D�ۙ��p9�<�a~aw��y�v$G}���14_R��5�!�LO��9<��3'͎���p.8�
���xM��]���b�5�B�<��C��Č��Ph�6�C�Ob�reM;��M�8��K��D��;q��M�'��0\��r�/�u��ξ�	P��1�����u~af]��fy��Ё bK@���h�%��uXq�JFy�m�,W礁 �׍j
"�D/�g�e�SH��W{�eD	N�ָv8��͒�Z������LN?���I	��^��u����|؎�0��0��a��ʓ�B_*ڂ��HM����1��IvD(J�0���mR�X�tn�}����eNsn��1�����r(����qT.����~��]��v�F������Uc/$��6�Tz�{tTP jm���+?���s��jTv�a�n�Y��q��%�HFNI8B.m��<8g�9��{��)��w@��s����G��S�R}�@���U���)��9�����$kK�Rr���E���i�6$�SP��s���l70칙`F[t������N��-i �����W�#D�l�c��;!��=�E�;�&"�w��z�r��q>�7S���0ek�p�ɴҌ�|���Y���N���� �Ч��!bT~�?��-�~�g�
}mr2�Ld��낰} wa���s����(��o+h�O!�s��צN�%��Nܚ&:s�s����4;E��&3�4��Hc�-n3��Npك� $E�ܢ	>�N<;r)�{���N�,ԡ�kO�7�7M�
XlxV65EB    fa00    2210�QƮ��sx:~˂��s6< F��S�r���Z�t��۞�C�.+��q4�[X���9�@���e]ڧ˗ �ޖꢁ'����*`Q�7m�.���iH��H �I�{o��z�ǌ~�o�w]Pi�o��)ǚK���x]�L���+[qp�vCOc�!p�`����?���J]�G���.~��	A��|�I����Y"d4��(���`=�F�w�j3��	諎�ؤ�Y$�/Zm2 ���R���a:XG�inc^���a�z�Ec��}�n��������M�,{�(m�,�w5�W�1?�@i�<��9�X`f�BI�k"Jޑ�WO��c�vY��q��j�Cm_�WPV�0��6H��H)Wg��ұOEv���O*�:��o���E�N��sY��`"��a._d�Ouh/��0�9���6C�0O�`1Ϙ��W �t���?�N�(�O�p�G�{9�W��!�f6�ݓ�O��%�y\B�]�H|�	�N�W��\������%�8p<�[ݽ�1�"�>Tͪ!���NE��$�w6�4,�x����˝�+�;����{���Ҏ��"�(@_ZMl��KZ��wmMH>֟c�eq0����_�������!��B�����w_(Y�Y}�)�8��R@2������6N
0`���qh���0�֩1.�	#�v��$n��x���[g�QoNɥ���y,Z7G�*����$�H��@�:E���������~�V�f�y����:�Q�����L�.�	��Lc,s(пv�.�d�SG�L$��ށZi}�VpRRk�m�����i۬�I��L�D��b��+�*� s?+�\��ѩ��9�o��РY*[�����A�}+�\j�?_��u&�>����D��f&wO�w�� S=�AjVn��&_��F�eH��hM��K�$�{��G檊���M��h;:`�R���\�y�tFlT������|s��Ѧz��6��e 1Ǘ�:����?Aey@���e���É"k*u��]~��V�����F�=�<X�̖)�&'�*G�T��_����
Wk� ��t͇�^�Ъ�;�����b�+���w�&�/�I2T&�aǴ7�7�su�����r�����`K�[1��y6�(���`��j�+�����S�bL�a�?wa�A�QX+�\�[ν2k��6�����ʷ���L��ai*mo(�{��~%���Ye�Ϳ1@:����2�*�u'L)Tr��1`�uW��h�����:��;2���e�O�ﶒFq:��(��Ir@V�s�s�&#{�!,pWn�F[:]�"��vϺ��0~�N��U��������ٮ��FT��Yǿ�_'��[	�*���En��J�M5_CVGS��x�Q�#��vB�Z(&%���p����2NꂬIeF,_�v���g˻F �UN�{�'V�2��q�:!�bL�����IS���?�=o{	�-�u[+I,t��M��UY��/a�Z�ON�!��2[d	�#�:.��]6�
�1O�Oˢ�0-1����Rm��̂}���>3�eK���B�ld#�s-p�1祮�y�;�W��ρ�F�$�a�i�Ս�Y¯�uN(��������nm��uq@.��Dc���|^�Qw��H��G��+�l�����9�=|�Xff��1��hNG5�n�+�y�G���'pY6;9������$�U��[�A~*	�D,ŒYp(��Q��1 Lo����S��^O���н�����|c�u��k��D�&IH�&חPނ�<�J�~-3 ���3C���OMξQ�����uma�}�~ y ������0gt��Ä��"��b�߀�>����-����~U��1��˛Ug�BoT�h<x}���_
��"��Ԅ���y�6���Ł�r	t�O���#ygE~��s>�����w�9Jaj��s�o��AB������6[��D�Ӑ��=��ګI���"�Q1����i�R~��^0!C���f�|n"�'���k�53�� Z<s��e��9m�&BAI�7Y�F6���P%�7�2�]',L���Xz�ౡ��ť��	 W�l�k�F����SG�B|��X���6��|m�ơİ�o��%P�M��=��R�(T�K`��]���`f;�t�3���G?X�'4g��8�!~@��o�D�!��5�(���Q�U�	���6oWt�c�ҡ�U����7�7��E�W� x��t�e�[��Sr��΅��Dby&
2�9�-����\�,�g�B�,k<��OUV�K\��7`���j�OK�t����y!�۳�X���65�=���+��'�(��zh9��>�q�¶|{\�P�����tSH�����^���� 8�̙ު�
�$P,��n\��_>�?��R(	����XG<���/H���GxfN;塿���5£p�}�wK�8B��TX`�ΐp���b�<R�B��	�
��4AP��(�	��e��N��A=�s~F�=w��f��ۍK���1�=��l�E�1������m�m��fE{g(����dm�~뼳L�lL��x(냝&������6ۣ兙��r�8蜬&q�m��ɰ�0x�0W%�8��������3����S�'Z�|A0�J<�s�m&6�]�'wL;�Xt[�5r\֭D�#�:��y�^����61.�g�x�jb��k,������`H	��vq��{����q�oz<:_��G�� S��V�`KA�C�I��om�D��i������T�/#�c��(L�	�SP'��')1�8Q(��F����s{��8/_>Dy��Np<�(T����DK�T�+�m"R��¶�<d��j�M���cP~uӴC��d��%�^�*"��pd�]�DP��N���,��	�j�,�4�[���f�����(қ�"��@;| �9��9,�4�ǶsQ��y����3<���n\ܕp�Vrv>a�R�or.�����B8�9�m��i":^�^e@��ɕ��2�����O��^�tσ۳OA������q�"��'�ah@�5��[�#�D����+�g>3��糰9�������ԧ��z!(}�y��5���yQq�r�q��	}g0���9������0j�Y�"Bow�������,�w2 �&M�x�X$N�,�w���l�Ѵ�?=:aԻ�#Q��W�r��Ֆ5�!�r�*���ʌ)lYI�5�?����=x�ɳ��ɦIr
O���?��vʪ͈�#�]����	��~���<�J�av��ky�qI���BA�����IĠ�~�FF�� C��<Ctg�Ռ2��ĩ.�8�{+M�.�&Q���?gӍdlR�� P�Tw7ϙG1�|ߐJ���J~�1��j�Sf'V��T ��W�H����X�ln"�;A�l(��$�%ڀ�;�T���Ť�[�N�?�*6u�1���/Q��� �
U_��^ HTƦS��s��ϑ������]�k ��ķu���P�^�ZCq��<t���GT��3�#ݼE��y�^���gR�Կq�З7d"�au1���2`+�Wr�:_����#�ܓ$�U,��pN�`|n q�O��Ծv�==5�p�����}���7$E��t����,e_��EO�w�&��x�eb<�#�S1����S).�e9ϰ~>� r&��+��;ÐEp���~�vRIh�����z��|�p�߉H5�p�q]}?���؝�V�2ɝA!h�y�Aݕ+Ύ��w�C�*������QX�_���gn��Ӷ]p\��`��K����y�B���IY�*1��-����\�q\�,�1�S:TGB�C���eC�V_�Y֕�qJYq>�֍p��3�Ւ���y����֭pR�X���3.�
��;���������V�G@��}+!g�.�9�¢���r39Z�ً7�(�X�S���vk��hFȋ��n$��R�n��}�,no{x`:��Jv�ο�KB�n�ሧ~ʀ�ɩ/�9���+;O��dF�ڊ����ʭ���Ap��mzW<}|���.�2o��dՙ�ҷ�K�NE�9���vL�����!�k:18#�yO�/��+�&�� ~ӻ� "n���9<�ڂ��M�-�J��?��:������.������=����2�	?��S�	��"[l���t�Ņ���؍�/�i	�L�v�VP��2������X��=�qrS��?�X�}�$�xr����z=�K�|�ݲ�C��S���d��da���9)����UZ�}j�/2��٭}���DQ���fP����-wk~L���Z�s�>g�*�o�Dd)h���ː<+ ����\E�q��ǟ�D�Z�$���!��Ɨ>��C��C��{g�4S�z��2>��P������8SO� '�_���T��{8cvà��+���Sa��ϡu��%�c�/�����F�����4)��Yə�4�3Gϲ�y�#�":S���/f��_�N\
���a�d���"!�� ��R�x	dow�E�� ����OX*~~W�3��Ex\U�]��Ə�QE/��Bg��m���?O�6�ws�C��/
�.�Tv F�3W�I4��&���'���)5bKک��D�[���;�n��S�P�F�\���{��;���=P�XشL|Jc|D��J0��Y6Co�e�$��+�huF��w��E�&xXBӑt�����E��_�u��"$�\����c}�ӖF��=��~�a�Y� A�:�Ǡ#�dS��]�ܠ���W����-Rrn��K�Ԧb!/��}������}��m0�aS��̍�~�_�*��g�@�TC�{�l��l)&��?�;�]���1�c��k�ᕆp%�((�Ŋ���Z�Ǐ���p��9�w+�eôAwcU����>��Z�.��j2����7��7�PNr�� ڍ�JQ��"Ib�lL���XL�a�)<��6c�_�h�Ƙ����2r��E4�;԰����٣h�*�r�	EW��������!3�5t��?g	����=,눠���*FaD� .�C�6���p��n��G��{�T\��u6r8е�9�k�1�D��1r�ti���d\��$����(]��v�����{�0� )5��d����l� x��"zP�(N_.�]#C���ܑ�	��k�����	Q�'��Oe�������I�펎a��`D�<�A�;�.��5��C��s�B��(;4���yt��6鿠7��;E�8?��T7�8��0��s�A���LR�t�먓�q�>kY ��\y�4�@��$p���F�0o.���G�
l�3Y�\N�[nD�ٙ,����\���Bq��.�t��B��,!a��#I6lhV!�(,̂lp�Ht�q*���,9*���*��g.�r�
^�w��w$6� ��"+S�]`J1ц0�ɞ��o8������B��^�7zP�cJ��Uu�9�g�pn1�IG�����)�
�g� ��r�G�Dj��h_]w�hS}v�[)Q�J�S�{P�i�g]<D�gi�_	�
�x��#o�V��b�ϗ?0s�Y@zt�*��Q��8�>V�ʲ���9R���V���4�dW��E�+��l����X��_�7U$�)aqz��G��pf�P0`�!C����Uj��G'�Q��?��� ����&����?x�u�!��Q"Xե����D9T�Jt�5CN�������
����B�����
c*|,_�N9W�>����S����uN������bE���]�|==^��pb�]&yJGpAԔ���1eR�,	�E�P7�40�H��S��7��N�wU��Q��6`PZl��qa&#�����l�0�֣��hi�X�$��z�(�f�q�7$�G������d|-PA���h[~�P�T���(�t���.�x	T�媅��GtQ���Er�^N�7e�&����B}��YpK|��@�_z��$+u�wU��읡ѥZ�KF�-����Ih]tfc���$,�;������A|~������o�C��o��6���x�E�Rn�+��w�������uiJm�IḰ��G�p�,퇀Ӛ��e�
��&�\��#G�Q�����q���C�U��:\5HRd�阋7��|?��Y|����r�
�Z�d��M>YZ�ĕCm�`��T��~���QY����A��p��9R#ei�_�/AN��,E��9�L�69���!����ͬ+�Ks���<L���.����:eoN��{�f�0�N: �+o���0�>�u�j�D����7��f�����U��Qh�*H�-��I&}�d�'N ��h���G`;�")v>J�}��Y��U��2:�:Z ��sN��g������hׯ���,Q����SQObW��0��~)��{���������9AQ߀�ʥq�#����R���y��Q����%r��ᜎ���'�=ljP6/g��(���BU�����TR��<��J�i�f�3<�1Z�$Rņ}�?���>�ה$�ǀb��\���?#5��ي�b�6ֹ�������g�H���|�I�yhH8���b��ˉbk&�R��WN��Wp������Μ�݃�+t.�{^������ʌ:C�&��{�_�yW�M˜*v��7�!���^��Ȱ�~�gd}kw��5�@��f�R����>�$�BVʠR/=�OG���4�L���>2��s��yvM?pYp��>@�xk����ʄ?<��һ#��D��0k�ϝ�,�5 !0���aou	�{�����;XB¿6��/�ǣ�s|?���*��������-��n)�i�@�r� a9ÌG��;Ѫ:�C���L�yzt-�M�23m"بrj��Q)'T��J������	�р�����$yFZ�g�X�8v�/��y���\�}��P��MR(%�GZ�놥��ǟ�6��g�\��R���C�?�^xsj@�%�'N�<�~'�_�Y���襰zU�xA/��oǳ*`ژ��0,#P�d��AO��o�H� ��f��V���d��ɏ�Iz�=���T�@�\R��Y�z�ep�)�R���Ґ�l�.J0��M�-�/��^	�OR� ��.���č�&;�9m1ϣ�"^�[��(&��'�ISK���?����{!��c���щ���%Gt��x�g��a�X���Π���/q�����
���Fh�1���>|6�H'_�fzƻ�{��V%�.�z����Z�������k&t����Ξ�Bm�NO�w��o��*�6��d,j��X0�mg]�̚�s�D�^
���c����,� W˙	��o�o]QE������K��ep��<G�'o����9B��V
�^�k�v>��'�k����Cu�);�m_�yxh}�&9ȉ <�a�|�+p�I���jU\�!�c��2��{3u��D=�cƙâ��pK+F};1Ο����}c���W:��P,�vp���o�Y�Ő��g W�+cB��U�@<.3�M��T�Mo];��]�U�x�
�,���D�Yv�
�Q�!
L��- �|A��j����ǎ)�
[�G�q�Y��Ndmϱ#z<��}�d�d�a�V�2B%���&oY�j[�Yo���*�����y�[�����`E��2j�����ZAUHӻ�[ ~�`ǵ�`l�ع�G������Bޓ����6�.������<�D4�(ogv*�l��&qGT�* �̢���l]wB�|����-FX�l���c�8"�T�S�>���������:�����%��g8�%c( vեUZ��Q��-�4��eu~R�%�b�(Do�כ/���I��8p��R���Z��fA79!���£��I2��&���M�D8x�w[N?	�ˊ=�ᗩ�yXӉa���)$Ju�ӽ���\v ]W|��Ed `{������3�=vUDw=[8yu�4v,�KcL�����A�<�G�H���A��{�Dа�2/)����Q(�����-�f�~nVHi{���6�N]��5��4m�:E��u��B�\�5{�JF�,��dg��آeg�Z�xXJ��+�e~�LVo�?|�+ ��)��`��f�-�b�d���eLr�ªy��QBE���9�K"�5�i�#h��m��m��O�R)��[�����dw�}X���<ފɨ��H�
(��O,�߄h�u��ѫ���ӊ�|~	�z�E�-��2�S2�N��_���"PSBQ3���Gi�(v5Y������P��.)����_e��`�ޥ4sT�����
����'m�tj�X����o�rN����V�`v�9Ee����L"�X�F��(a�ƶ��TP�h09A��NL�6���6�]?ﻓ[�C�?	�����&&-�=����6؇���F��� �y	Xal�����og
qF7~km���r;�t���*z��U��&����^�%��2����_D�����u��,C�D˵,���1xr�WZ}�6�m������]�\���IT��
5_����./�(�Þ��6���	{F0և����
7l��f����f=(�����b(T+XlxV65EB    b396    1ba0m���*w+��DE뼢���p�:g���a�wǂ�;~V\��gGePr*Y�Gv_�_�s�j�v]�Z� �0�߶��dZ=��A�!�n6�:KA��!����Z��b��N�,|��Yrr��n>ʹ����S�{��?t��HM:��p���;u�x���	M��m�%�V�r�e�Pm2��c�/�s�^4���>��W�[ ���?E+$��e"?�l��:����V"'��<�1=���^\���:Ʌ�(��\%���xJ���v�Qc]�U����7������Ǟ��q�laI���q���,����J��m�g���jE7��������s}�� �,��Zy�D�dx�1��`��	��"�������/o��pT�c�-ϻ�pk��@�d�\�@���|��7}HMu>0#7W튣���!Q� �G�S,~��\gN�	��Xd�x��Vm���Y�0���^�_�ͅ�s�9CFN�<&-�h�ΰ]���ܞW�)O�  ��BA��=�a��R�(9�6���K��i���	���c�
��+Jl���m/���Zq];l*�B
t���� C=���I6�SQ-�Ť�W� ����G�]��uI���3I��ha䗴��<bp�)@��kg�}_$0s�+�.W�6М�M��[���U>q&�ij:PN�(ȃ���}�����?�Q���V2�=����`!�T�x.Y
8�c� �����u��<��j�L�����&7H�u%cӄ�`I;�#���ECZ�ѷBb�v@�p�Ú��[�we�#�&HJ7�(�]C\h0׾�EW�����w�;�����co�X�5f�y�/x��������c�$�Œh��fB�q�f*u��#��z"y�ޭ=��밾+��P�9���E��'nufM�/�;[ ���髉�2�H��i�z0�}���y����e��{i��/�*h�g`�B�d�Y�M�,������(��Z��Tm�"��Z��t��1� ��ڭ��vT�]V���v<@[e���	w���A���`��b��=������*�/�x1Dz���=��&��ų��8�!�6(\t^��v���m�U�/�C)�������̻������ǟa[V�H�=b�F	���fHT/�B�hΆԕ,ݙ%��b���~ɣ�����4���t�RS�+�H���+Ƭs��i�t#���p�A�iU�wXh���~I8���:C�O�\�=Eah��<�?%�D�tPjX���o�i!�L���e�������+��(�%D�,�����_4��;����B�A�f�%��a_*79�ۅ��$zv��1�х:�': ���-v��]�KY+�(�X�\6ƹ�c�à�Ж{���pj���hL��~J���Dͯ��Rdp0��\m�}��?|�:S�O�㢣������z�͊7Ր�!=�)w7���$�S�(��/����mm.t'��Ʋ�yUZv_la[T�S����<ƒ�C�����3���:z�]I������U��U� "��D,�Ȓ2��B1B��}N%�{{�<�1�����s�Ngpd�0ʽ0EpZ��sݼ˝DrҌ�=\�/M��#3� �"Şyn�s��O��&��r�n|K�z�%�T/B������~�~�Oqz�Uo�;��r�c�����F�R,��K��ð�C	��E�W|��±1�r;3*�Ѿ}��E�-�k�	���w�#�BE9�U�Q��8̣���t@BE����y'%�ׁƝ����WL�Ae�|�Y$x��m������5W��:u!f��f�������B�AJ���e�Y	R.��H2�&wZ��0}y��pT8s�4�ꍀ��9����Q�3�!TAFF�jӃBt����%D��-I��7�S�(�F�DQɹf8 k���34�EN��"����X�	���q~��c������?q<*'��$E%p��E,���y>Պ���c�:�c�m�ܝ��%�ǫ��|� �+�o�����K�������L�v�L�]�g=��.�B�	a�� �>�I�:�C��YJ�O߫S�� �o���Vz�����g.ʶ�	k������f@ �Y��?=<�O�U��}	q�'`E�������7n��a��HGV�jܑ��wf�&N�	݆]G�E<���3*F���<%K�Ȏ�\�b)�~��2�ʖC�ֵ��N��a�M[�Bw՟AZ� � �ٔo9�Ģԫh=9��5j��$��-�����uq��Y����Qqx�vs��Б��f�YyBukD��|P�����Z>��=�l!��E�\ ���3��)F￮��pb�]����W�,�B�ħ� ��
uX�`RW������(���?G�� ����wU�K�y<�L�܀��l��:�
���/U����ep>����Ǹm>"��%'��i�N�8��E�]�T)p�/�S��H�M襁[wE#3K݊�ݨ~S�d�k6%8'�O"�!�Sl�uF�6��G�XU37���k���ᠽ�nl�����'���O���v�:�+P�id�O"�}d�/j��� ��N흮�nr@����"&blQ'5+��V?ܖp���bK;����� ��{�p=q��	z,�4�Hy|)��ǧT�	.| |M���#o�˥G7rv<(���;��H������6�{yxGJw���=�K�T��x�c�%8��d`X��?v��gP��z%�Y�F�<�.�b����[�D�8ě�����K��Y+�^��}�[r�̍�y̲+��ֻW�3�v�����wu7�1 �o_��|Y7���we�)��GD��8�+���d�0L����[3���t���U��.�{��[{AkJ}-o��,�1����Ј:�"�؎�̛b���f:1�yj� �����7(��|Ϥg��r�\?�;#k^1M��o��-�7��ԫ�滻�Ko]6С�:�]��O��\�>��~�|:/�ep����ש~�:����Kj]��y�w�=��޻yr��@�u����gV�b�@V�t�#HtI|�H��;�%�_j���P\�{��w
��7���(2���1X{��J��u.��b�ש��Şw	��y'���|�1 �{��=5(�UVla��^<f�Q�u��\�z&&y.X-
x�$��E�%�g�k��&8j���X��Jnd���M���q4N������j��OY.��T���bc!��'��"!0[/]��b-Q�`i����;�z�{�P���ҳϰ!V��t��{M[��b٬=�lg_s��-6V�qqnu�`�e^m�[���Y7d-�9�K�Bs�7��"��E� JL7��i�G��^��b����Y+�Z��� r'،��ȟ�r����;���e�/E�b
)BG�ԥ����L�*�Q-A,ŷ�+dp��vJ��A��:S���%t�����ak��<~�#���︨�cy#f
x5��>|e�,�_U�;qqo26aS��CBO�h��4�V)�e�Y�W�.�oȚ��H;
@�2����}ǁ�c�B� NƸd��#�f�o 	����V�xU��U}h�-j��=(9\_������tiF������d4��M��Ź�����������-�[�9�޿����m��Oa�D������X�E��FH#stQ���
|��Q
Ⱥ��j�R۽p>���2u���|;6i���k�=O(�c���yK�^�Y���F���˻�~�b�.,ui9�ʱ*o���� 3�>/H��]��=u��(x���ŏ�z�Ҕ����!\�2�ΤS\���kΨ�*8+t��#c��^�>	��iX)K��LK��/)n�� �f�q�xR@��N)M�\3V��TR� |:�߸Fe>KC�nwpD9yJ��{�x��tSG�Q�ʕ���m_ʱY�u!B�v�k�C�O��fi�>+Ql�W_����lk��z���3<��}5~t��R�g�dv'l�ŪB��E8��|�:�����kt�c��6��Kn�l��[K�$TI���Y9�������n ��h1ܱ��A���2�>�b	y�# H9�F�g�w8h?�(:���+�)�����~��s��-ўMWt �X4=��U=L5�/���f��=���Fܡ3ao�˿W3&��=��CV��5�w8���W��Б%:��4��s��4=���( ���# ��{a�<Ōw�����F����g7�	��ih�"ÿo���.$w�i�[�pyo��Ac�Qcm�iq���Վ�9��;Z�
��K�^)��;"#KA�YV :�꣼���K$ܺLX"g-dE��Dq[.	���ј���a��!\ ����}���L9v�c�G��)��r���3b�Bا��S�Bd�+p1gkװ��{
@;Dd���0�5�{v|h� jO,���}ui�nH�����rA�|�)<M���?g�������&ȝY-mJ܇�cѐ�ES���{������ڧ�f�pMqu�\k�iQ?����'cn����u��Ajy�����6RQI�H�_�DS�5��,rM2��0�C���gH�xZſ�f ���
="���iu�k����B�
6��ӜB��6W����/���ϷG�&����|m �U�j.f_�0�\�:��^[��A���H�h��O�Ȃ�S!ewR(u��7���8�b`!6]�Ӵdph+ͱvo;nVK���I`��X�����?hx����4"+�p)�E��r6�R�pn�}������2��8��1���Sz�a��!⁤�5�.����ʌ���zq�c�W3�>�n��GF��H�}d����XB���	�X3!θp�Q��K��š���	$�4�n��;9[j�e����Jm
�������`n\����X*��I����y���.[��ar2x*q��2'�0��GN]���wL0D-yV�l�@�6�������n��˂�
"�8N1��!�_fc��79��<��H��Ƹ��Fh�o���7�B���9�}�k�x嬆<�p���s���]y���v!��8Q��C>�����1�6WFIs�L
�q�N1��C7Z�9��A��G�`'w��Yt�g|x�;Ys6��Ϩ����2,JED��L���ɧ�]��^q�p�b`	�:�G�3I�;!ED.���I�·',�����fQu�TW�dJ��Mv�,q��[l ܟXj��{Ų�h�w��0E|N=��U��@1��|];��w�r����zf+�f��Iċ���0H�0�T�r(��Ƌ]t���B;�U$zF�xlW�$OF��)�!���.�q������'��+����䝫��Eo�0G�tD�i���Ёy���*(+���nP�4|r��5K���XJ�N���{��R/�F��7�g�pʢ!�ʡ:C�T��ؓ���w$t
~{���U+h��=P�T~d(:$-����n@�"X��t�֑���A�Lk3��qj\�;=\�/X���F���D�@�i~F"���s�ei=P�} �O�����p|.� qR�-���T�VA�A2��_�*37�n�p]�o��F-]����1��t�d.�eȤ�>�Z�H%fo{B���4V�M�#�]��?��%!J</�a��:����0���b���d8���g�_8�?XI1]"�̯�������ZW�no�.v1�W��b����I�c�l
2	�"?P,H�q��c^T�A�cBSԱ��j�N�Z���v;��,"&���ȴ��Fn��k��3g;f�!��6T	G8ڄl���ru�<+���2�鲭�.ϩ[�>�� :;,��u(R;:���C�� X+w�"b���mw�teIm�	�C�Oo��y>�'��0H��j`�%��T}p@�e	�p��dޏ�uݎ��-i��c�u�����)���́Q'����Su���g�f�7��-l�>I�dtݦ�d~�՘0�:,�JV 8F��H�󐑨�$|�k3:�k�Ժ�.��U;[����R#!���R���O�B{��Z��	8|����P�nY��Z���+�1X�ކ���։��"�S�)�F����Q���h��KiS�J��� �6��1L�SvŨ�}tɪ����uB��[���@AH>_ϧ�!P'k�X?�2I�q��$�Qz2=�G���ɝ���Pϵ�Le�AA���0ƥo�`2��IK�D��P g����4��:�jAY�#�\ӹ���/���,x��������Xb6�;��=u�!�Ċx
K�\�o��J2����'�bH�q�t�0N�~�w�-�#�8�8�쥑D��MV�4 z��.x.����5@0K�ҁc�`�כO@qcI�6�׵�S�Zs��c97�� �G.��l�U�����L���/|�O�>��f��g�;��>J#������������3#�JmZ�%�e�E�����]���Of)6� �Z�|�|8M�a�
	�x�R(���f���Q�00�G5%�ʚ~5�Z�H��W��|U:�H��H��xy�l>�c(Z�-�i�r�NE��HU"�5��# � �NK�j�6[��}cU�JLH#r�!�Ϝ���"~�.�ʞDٷ�W����*��K͘�8\���]*gM Yl!ҨT��c���^A)��� ��]�'�w|9���
8z���i*j�ag�k���ίoBɪ������bk��c���fL��YG?�v��w��s-��P �`�o[�Sl���-{��b���|o]�Ռ{�rΟ��D=V@�$'�
T�a�<6����,��k�?B�������"��y��?�ѐ/j��7���%�H�4�P��]�K��ktr��5�������_ �f���?D>�
%Ӛ`�����g�C����j�u�$�4#�����y�:�����f�5���صJ[�oz��3��y����2׺5&��a(������2`�R?d5���괍O�[e_l�3j
@/�JN�����1��[
��N��i=S
x5b�|��pV��aVM�e/K4ݮ ����
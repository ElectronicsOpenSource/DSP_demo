XlxV65EB    b060    2030�,A�Bd�.���m]�vǳ\��$���j�C#A���&����-|���_/J�}�%�-���C�C�ʹ�?��q�P~�Jh4z��)�ϫ�w�d��XP1�L�y�h�N����QX uF��HjM�s�$�N�؀v�D�������U,0�5�Qx�i
gI��4�n�+�}��$���$���SH\9o�~��u옅�5��
)M�����g�1RvS�]��&�����ߌ ���	�*̼�[ߋf!����������+�Ŧ2�4i��� '!�'�pR��%y4�qE�ȡ�.{u%��|��y^%���v�i̍%
�8+'e"����j�#-SA�2G�xf\�M��aB|#E�R\S5k�n������:��
���ᮇ������t�!*�q]�q�mUL���-3.1�b�-�xnф>�+�(4Yn�i.݄ �f����hk [I\���x����� �<�_�ahN9z6/rR|ɸm5��h-�ņ�FƟ2�����;�j�;E�m��ǝ�C��X����Lu4�T/_1W{0�`Ku P�ɛ�ȁ����vb1�x�7��iS�-��i��Ul���m/fq׸R�U
�ht�v/S��iaI5w ��Z�$N�y»l�۟�₣��M�:��_m�9��5w���ߣa��ګ�I��bs(L� �k�>���5����L����c�٠X��8�,04e�?1@��O���ӗwVt��
�
X�4�@G˵s�z* 4$����7Z��G�ݾg��&�m���2��Չ�.�����?����kꘫB��=��r>h/ �	��ݓ�ػpu����"�%n�UT��)?_A,���V�-وk��w\�9�t�!����2�b��rm�嵖�yJ^�/�oM)�>�"W�*E��[��H���h��k<��rr�}
�HZJ<�eɽ�L�	�}�`����ұ���ѢlrƗ�Wsiu���|'�Y��������:z�,�9Q����pMcz�.ʟl �p^rL��H��_��}�4�y0���o-��ϻ�k8�����^q>��Oݝ�_v|
�ʟQ��S�/���=AIV~f�Oi������"��7�KX�����J%XAa�����&w'Sa�!dߡF�6��A�Y;�H)��~�K�3�\�[TS�P�#�V̐�v�p�.
�vq�Kj#��\�ɎΖ!x�k�Q#���lHJ,R�_g����*M���-Xd�a�<��z�+�L�d�d�z�������n�נ4��j�D���J��\ 0�*8��-I��0��H¥YKh����~�F�P��`����k���AW�{uY�Y�)ז�����N���4�+�r۸b�׀�vsVW�ɜ��֖w������R(�I~@��gL��������ᚼ7π�9C�B���121(!���?_s���΀�F}����/�I��]��� �:��e���A��������ޝ%�$�}r�R��z��[W�6������P8�G��<�^�0̖l1��~s)�}�:�0R�� �i�T����>c3WC0
�8^U�:x������5FAۥ��%��4���{����M�l�Q٥���4��P?e�b�е���a5���f_�#F�7n��-��nR��N�$��R��,����Ȳ�Ļ��A�q^����Ei���g�� Ƨ�2��z����=q�L��p�蚟.�5�eI's���Ψ 87g�n&�))R�᠁�k�2�I^:�O,_�P����v*�5{�?��c5�?v
�o:���n�0��Z��OuKHv���(�����̿<L䊐�4AYj3V`��$	ƚk~u�!�X��HW����	0e\jw��柺3w�{����t�d&_c���R�[̆*J>�Lc���˙d���r
���2���F�������`�\]���1�[�#^e>�BH����n��No0js&8+�	�WF[r/���sS��qu�[r��&�o�o��d�����G��n���갪�`��σwr�I<5�|�^vIO0�4fb�>$���BPWY�i��a�!mM�'�sa�ΐs.���I7�xK����`S�\�f�m�|��g�VlNsܻ�h���=#AЍaC`tR_Ζ.Z�N��k$-ZՂ��� N��������R�Vz��Ю�4�L#�9ϑ��K�i74eAװ��޳��v��C�j���h'��.M~kv����TeP!T�;|�`��|x�j.!�����L��LAM�_��bri�����ÓOqF�-f%�����2zmؤ�+���m���l��V�]>�Z�i�E�ap3�)%�.ץXgq!a�5PcNȕF�^g�f��'v��c2�V�#�ߙ����}�9��[���C�T7�f���|e�����e�J�.h;���KLkt:�W�31k�.����!]Ѩ���䠔t���������E8��������:-b�Ae����?4*=�B"J<ػ�τ����j|�Q]�:�N��jrxȆ��@��;�������)��v|����I������Y�A��U���{K������7�o'@{�����>]Tf��:�ݪ����q��S�����t"��k��߃��jr>pF��C�W���������T�&3��QAx'bV�e�ˍ?��d��qK)Z3 qc]@ɫ�����Q���\L�O��fE��$��xO�V	�x������v���dC�d�xt��EHl��o�h�^D,�ڭE�����erE�L��c&;)��.G���6��&����Kl"�������5�m�k��W�5��^~8pE�u	c����Q*����ΪÍjC��8�.h{e����皳f�˖��P7<�t��a�עW|)�{���PG�Ǳ,O}���Lg�RIIƸ�\�).C�`kukZ�Cg�x����P�f�?�K+�G�7`����x#��aC������|S��I`�G�[8��N�>����T!�X�D�*,��GsN�������[k��b��C���]\�{7�u�K��ނ�=���G^�Ԉ0��6V����I>�B��?j\�`��11 ��"!���>&;[c��t�밬��~	��΅.�^�m�d��(�)cQ��r�ؖĆ/m�@�D���A���kιm�Z�X���ߌܚ~9|��3Y�@��㖌��.�����c��A�;+��A(F����i,Y���� L�9[Z�~��f�,G|Db�k�%n~�u�\�3��u�ߞ���D�tggĪCy:��͈�#N��v�lQ�#�)f'��n"���m�@K��+,�O�깗&?l>�:� %륷E�t�X�4_� 5쥤c -ղ�i�8S�2z�u,>d���b����h���	��r.�>wX��w��6.���4j�D4���r �i�N go����-�m`�LU�w�P^Nm���& b�-�`���7v��fN���
��)&��,�f�M�ݨon�!$����������r,�[�l7�۔x?�����K��2OD�aT���bu���5YM���R�r���ޮT;��C�<�諿�xrk��~P��� "��U�a��<�ɳM�Ar��7Bs����1{��.�R���v�P]�f�R����"B5g]�����6�+4�4fܺ����&�/�ŉ[>��Nn*�"�����L����=�) r��奫b�Y�^�΍w~��j��2C��$���P�J��Ů��������l����!�F%� �h�m��H���Zpgt�]N�.m��M0!tT���QJ0$.t���xF����0�q&˥9���6����c��] �?'�|�����=�Y����:8�љ�U��p�ܣ[y{гCLn_���I/��> ��*�S���]&\���֓�2�oy�C��}���5qw���9Y�9��L��d����ϱ��G�bc���h�ϯR��H4��3DZE��i$]'tp�Q���z��|Q���;s�&��F
�
��|Q|�0Fn��,R��C��ܔPBd��}ةZond��rH���w�Q�qTþkg	̚�tZ
n��̭"],(ި���G/�w�V������A6�D�c�t����#��������O�f�<j$�l�Y�WO������~q����-F��w�e���]5`��JO�l6�G�W��#���5?H���Z�k`�	]���<��}�In���m�g�� �BE�K&B�:���.Yʤ�gl�j�9 �ؐ&ԫ_6�>}��"�^1�tۡIX5���c@�/���*���CV�Է���4�Q�A�*�������3k7N-Q��K��-��:&���H����W�g�����cU� �S0�5����5�dŠXM}
PFO�X�d�z��X}P�w�@[C:�-�Í��m�D������_���q:5�d���*�.*�EY߮��n�����0c��T���0dݤ^�g�N�Xf�v�m@��re.3�@D�\���p��R�?��������������&i����<��l�X܂����T �Sn���	���B}�K`�s��a^�B�=@�{-ބO�ןlPT�ݝƄR��|�R^�C�,�^K��z�1Y���"�r	e���8E3��Ǆo�Ӄr�lFx�|��1��F�h��=%��-F��h�ۭhGA���$�djQ/}��$a�c�J���l�&��Ϻ�U��@�`��w �Ǘ\۟J=���Q�I���.���Mx�\�Bx�:�9<x�8�P�+��˅����#I�<�w��<���}f�컏g:��� ������9��+������8�DY���k",�}�4Bp�׶�o���P������;A��-v���/���i��W��{��2�Vu�y�_�>�D����2P3
��n3i���n�D�x�B��l�k�H)ȩKL���^g,��������ǧ*�X��H�-i_!�oE�Q�axV|Dg���mL��8��?a1��;^9Q�M�ź���с�DqmM�S5��Ғ���o�'�u����&$[��1oP��T��{��,&� �$�l! �Q~���\>!>�OD��8!"�Gc8y�L��J��R��p��C��ݳ��ck��a0
����5�|�#'�LX��ڔ	F�}��-cw=^�8ܑ�&��>oZ4�Q���ٟ�#�
��O7S�Ϧ����c���!��h"���"��
��L����U
���s���xk!��ſjP��1R��'�	gd�}b�
YA�d���r޺HT(W<��=�2��fT���s�	X�o~&��qӆ���Ԥuo��Di���a���R�jS|�_j,�7=����S������I����
RmC ��%�AܺR�PbBa�)ے'��t���������Y��c��bOE{��� ��=&iw����,:��Y�oW�X4�?R�_v�*=�};B춶�0%������vOtܫ�����YG���W"��-W���ʵ���.���ڲ���dY�q�7�i5?�C�L�nV��S�Xt.pvt���ʙ"L�����4�n"(:`�zJ� 1�y����N�.�,�˒��s�Ԏ���cǪs��W�;��<��j�#,��#�|�v}!��4�5=�!՝���T�UiݻK�7`�@Qƹ�H�����w��k:���d����M��r��j�lw���	��7�r��
���������AD�
ҧi��U_g��m�Ҋʗæf|	���W��#c�U&�)�Cxe���}�Бv��U'��VVJ*��D��aM�y|���N�X�lwq*�Lh�"_����{$��5Xf���i�Ϩߤ#@ ��-�����~L)�/T�sN`��8wK�� ��"EV��ā� Ge�"C]f�$�J_�PW�D�U��z����g��$��3��R�Ɲg��.�)m�t��]A�w��ɢ�Q ׆K�w�C��M�[ÆmJ5N��QX��X>j��/��n8�{BK����/��9CU_!!t���M�߫*���c]]c~�����:���I$��S�-�����9�юpR�?�P����R��ˆ�v����%�\e�f|��.@�{���T�6�g��X�?ã�nz����P�=pu�q��h�L����u_�{Ӝ��HbdN�N�L�Sˢb�f;�a}=�p)�b`�1��7)!Q\�n�nr��+̰���RH�b?կٛ�P�g����଎��$cCE�U��n�>`YJ�XF��&�����Xī326�F�=�u1��NFM�^�\�@�&D��TߏR(Z�Q�s�:�����k��Uu;Z�/z>9#��ҙT��?+�W�m/�6��[����6m��5M�p�/@�;U�}�x����z0�8����d���=Q��Vr"�q =	%� �;Y�����
U���$���m�Y�J�ʲ�� �:?d��Ա��&p}�a��-N�ίn:�� !��ye�.H��>z�,4����FY�c�;k�kV� h~����Z�d����s��lV��x���P��:��w88��`�fS��@k��{e��3�6���dl�Wn:��D�8=���F�X�~5�gO��t�}�[
v�@z��U����C���T�������Ɋ�)`�\d]T�HLGR�n��Ud%j��]�Fn��U���]������`Z/�}	�3�*5B[�S�����6K�`�VeF�r�����O�HpLQb��[���S�d���R��HG$���U�uZNsNq}#���`J�8�>���;�|�
��ZC�"��W	J`�gt�"P{�a�U�u�{�����%ݟ������.�|˝F�!{ӽ��.ݱRj�A��F���Z좿��T���^�B�ѿ1G�ɔ�!J���iS��?{�l����n�67����+�֞�[@�%��)��V�m+�H�D�qB�Ą�c�=.���k�hç:��'O������>T%M��[tS�e��S�(�&+�����!�%k!0e[KgtIu n��q� Μ������gĳB��c �}���񗱽oX��S�%�"g^��$�����9Ѹ0Q�k�H	�!m�ɝ�AmP��+�$����̬�M�>u˙h�tW!'ą�����S-�И�yҡV�g�����[tF@�ARp���[�å�2�F�v:�[Ŵ��M���T�۬5W!vC��!��cTk'���}j��wr�,��qI��S�T�ʍ�%��Ÿu^�N�n�S��40ߠ�s��O������l���<�濂@3=	!���Wƶ�	i�4Zޖ�0\�n˦�=&:e�z��	��R����;�����ps��5&l�xM���/�I�9�Nq��ە>,���b�� 4��R�"´��KrY���6V^U]�w2~r��?o�=�����^��[[��^�7؛"]�o�Ql�f5
x�)X���Zmi���ד��N}��(���L[uӏ�!~�64JsҨ:���m �g��۾B��2��L#s�)�S��8��?��<a6	gR�9N0�Ҋ#3�?'g�]zL)����#�<�L��G�6]vg ud��q�?+�F�w1���|��]W�ۃu�A'�t���G����z��֠u���˒�Y}�v5���"松�QX6D�b΄�r�s8�ʧp��AW��.{����昳��k.�k�����H1+�8N���f-Mg��O,�I���f4�(B���5�6�|���Q�t�S^�$:�ťw{�$�)0}���_���xŔp� ��	��\�qO�x���F̪�}�& V�K2���^�w����ک�Ʒ/�S�Ǌ�:+�ȧn*P�z^t�=;mY�i�W��ә���e[s
��Ac�x��V��%�D�z-Y�!��P5���_�½�'���$Y\�9B2�Ե$�E9�Q�q��[�u׈$�P�q��ӰM��xx��t�6���I%~G4��X~{�a��HN;0���͇`�J"C���?����*� ��L��!]~��B��SI�	�˛_�[tUo]Yi�Rn��.��` ��j��y�q���D�r�
��BE	�5�3���aC Ø#�r%���Z���Tk-����0}[����y���h
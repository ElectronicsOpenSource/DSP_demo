XlxV65EB    fa00    2e50��A�x`���P�)eXӚ�Y��/����n���'pI�G��X�o	���r��c�k��%�g8/aq�yF�{X�F>Lh�r$1�F������(�������́ui)�"/���Z�D�Jz]?n��L�c����MDJ��6A��6�j�UZc�ȹT7EzU%���6�re��Z��sj�����*k $QƍI�L�o���.����i�喁N�r�:>K�YT���7�Ml�jϟ�{�����`�Z;{��S�3��\#~�Y�!5��p���+�S��4
4�O��n��~�f��-)J�G��К�w������D��"^a�<��c��!�5�}�7z�įӂ4�e̨���~2�O���X�
2�����T��0�/;K⮵I�����K�4�ܨ
Ꮈ��1C3��q"���A��j���jQLx�Ve$�����Jo���/R;'�7�b�g��8���<g���e��4�j�߉�9����ԧ3�����'�A��G��Y�!��'�-���^���I[��>��u�H5�U��鯓��NfI�pT��id)��I�΄/߄�
���k�}({��l���S��Ơ�f��������.���׉$S����"�	hR�9�l'߁_���TT-�lD>S�F�^�� AC�B�.:�Y�-?�8%�N=o��$�0;�d�*����X��Y�;?.mRP��t��!'Ł�"K��tZ�8�-�>1i�IG��G��2��:.�M�"��=Qg�j�T��5�p�̇wRaO~����ލW�c�qAF+<{9��<�m����O*�a��A��]�FW���ys#�C��D�{?��'t4��@��c}>2Dp䀎������Z<���[�A����H3�5fj[�oE�ٺ}0@�Q�k����!�a��E\v_�P��X���=n���]�1��r�G�R\�O`+�g�\}�&�;��Ɖg��V��x���%6U����;@�b�4yN��w���B�$�dtyyέţ��qf$�}���n�dJZI¿o���p��
�fD��}C�N`�6��B-	�F�)z�H&s7����)hƇ�'U�8
��@��(�ݑ�꒍2�^^���g��q�o�:����tw�|���ס��/���!�9�Q�.��B�X�b_��_����<��?��_�ߥq�l�� �g`d�EN,b�<�G-����5D19>aV<��£rg
�u�3I2�)��A$ס��~���fP{�y����u��a�a�5
�"�ߋ�;J"�dx�FI�|��*<����F�=��GD]n�A�����P���i�Mb�>�Cr���6�q�����F�Y�A�y�&P[>,�D7I��M�d�+|  ������͹3�S1�8b]q��n�~)�������@���(���nY���-�Z*G�+H�acH�s���W(��[�����X�I������y������G��ֶ�Z���0��M�5�ɹ{%V���p�9hN������R���Iy')�Pʤ�w�-��g%�o(��4��C��`5R ������~N"������i	W�������ٺv�,XW]H]��:{^�(1��!��7FNj�.9�aJz#[1
z��Rv?��s�ʻ��u�M�����u],���mGwP�琺a���M7~;�)�؀����Αɮ�4�ݸ��uVD.+���%�KР�U�>�r�W�X�
z�\?�dె��U��%x C���y[d`���Ȩ�2'P�ȸ���&��`�Y*�5{+ۭ=�*鱲��o��@�¿�e�G��_��Jw�&Z�bd�KhA�^G���3�����njA�\$L����2C�t��	p9����ua���c�q��ؖ@�S$�B\�'ΟT9)����ol�Cƙ>|�AOM y�2�]�o��Զڲ96�Y�6Ŀ��kI�C��D��[�C7O1�X\�Ʋ�KG�̂.�͠�:�F&y�����V���ۭ	�-�wqv؇TA�	��+.�����"Ǹk7X|ݕq��ԭQG�q8�Tz?����Es|'�W�����������-�&�ēq�/��	�<���`��y�3_�%)�_=�hX��հCJ
��7�Y���lD��|�^2��N/5f����6�,��={�q�a�"EǭA�P�Yrn��=n.E�tP�=���Q��-�)#�8��?� �Y�d�/�/т���d����A���eI�O�~^�?oqt��j!���� P ����Z��
���Y���6�����k��:�d�]TCE�)�K��k<� ��<On�Se �fB*��>���U�L���
����_P~=�DxM�/P��60/���X�����
ZT`�U(&s��b��p@�,�(zS `�ڮ�2u�ӃU���	&��uH���Ç,Y�+6�_����a>�͈ɹ$ԮNq+x���\Ǆ��<<B����?��ր�]mhp��w�}��$�2&�؀l�D���%F�4�h�l��M+�ѻ�ML���������Yn^�����_���C�R��u��9w"�U�X}��]s��<3�٘˰PM���[��e�v�ı%rş��M�@ok�I;���TK�.�ɛC\��L�C���^�Iv����rH	��l>گd��3R�y���A^��	?U�jW��l�Nd���~?ᴙ�!04Q�2�'dV)��:iq.���[A�l7�钠9,
���ҍC��z��I���,w���Rf�	�r����Y��@&�>��H�ڤ��*���O�B����q�4�|sUj��Հ�;,�A�s�Z���.`���r��Z�w�R�,Z�6�"��%R«�K,���l|%�E^7��/j����}B�bs[*X�� 7�&��q��g��6��f4�;k+��g�˙܎��+!F�3)�~�r{��&3~w�����vW����8NG1W����7���z�'k
�uO]�=�[/���E�����@���:?@i����Jg��Bݒ[;�vӮ"HTZ���!�ƞ�攆�\l��'Bl�p�(��H{ɖY�S��dZ�^�*�.7r\i�/��\V�`��~�{9�Q�[���K���޺�c_�C�Q�j�����qo���(�k֧8�8R���=ת.v=��i�TE+��}����{pj��ݛ�V�!�pصgL
]�5] ~����X�=�Kڀ�O����`؅aR�Eg9_#}z;B%�I�_���w��n���h�}��X0 ����I��8��P��"�7ڇ�z�����:pzZ�ar*�����m?:�\`@���w�����N(z���X�rBXe3{��-�=o��K�RȈ)UA�H���jO-F����;H&��@�0Q�L�=�^�(§�(c�?��Mb���6n*yt�C�&'�������?�6�9���'�������A$�n�hY�
�ݹ -��N_��#Ȧ�}���Ǥ�/䓋�����o�O��0U����k�T ��f���}���=�H٭�	E�#���d;���o�H�Ji�(W��QfG��>��Q�#����Y��x�R�aB;rw�1�iL�``����R�7��G�/�����ϸYoJ��9��vr:!��*G"�
%�ϲ@����%��N�ӊ�6:Tǰ��3k�q8\�Y�U��9��s>��#C�<ԏU�e= ?����ّ8���d��z�tGߢN��q.��-8�fpyg��-v����!*�g泀�rԂ&*"7���7�]�V4�.��(�0,w���̱[�hmɥ�o�B�1���~� �% b]�))�P�)���v��T�aJ��Y5�N����w��e-���;I�%���e9M�}�D[�I?�'
��B�7�,�0�$�"��[/�T/�1u���i�u��|)9x�C4�qu������7�#/�`��)h�Y��Ȇ��:P��x�jy� ��H�_S-�R"���x-��n��(X,b�0[��&�&��)'Y�Ѽ�uR��ܒF��_���A��uw�أ��7f��QnR�dw���;��oHV��w{}3&$�.��n�-�'�'�TT�`[G��B�Rs��Yd&AJ\�sS�?x��{����4��X�ϕ�rJ_8ϴ���a"�E�T}��4�i���Q�S���F�!2��[��
L�E�+�r�2���#�dy��E�o��Ĵ[�G{7�ͧ9�~<���d����F~��� �^� m�:ފ��ŕ+vƟ�||ic��U#�<��Ho�4t*�A!f�mm�����І
�_o��pOQ0/
3X�k��
6WY�!���V���Ԋ����g�Q���;�M788��Ir�.�s1�ZӠθRa��k����5�j���Q\QW
��
@��>��{��:��q�ׄ����P*��������|QGA�:����>J)�W0�"5V��j�b��^��!"���x��ȑ�8�C�Ǟ�I�H����v�|U%�ڎ�d	���37_�f��	A�#������\��8:A$�7�Ix �sSD�����Gp>�C�/R ����@�"�_��R�N��U�Z��5��m��)�N;��*���i7B��BF5k,��B3���T�@���
�,�Q_r	͐�;S�*���{S'Ƿ�x�ӯ?ˊy��1-Z�"��/�����KQ�7�b�z^�P���*t�3@uL*^\���Xv���P+�q�g�>��:�&B;�Hxᕙ\�]˳�����}�ҙF��d<h3:`' ��^\@������vj��y�R`�S�:�SBAw���\9�ޒ�����)"�����6�X`�h(*uT�U
,��F��
)I��Q	c%��>WV�ۘ�|��ǟ?N<�+I� �����ʑM�A��6���n3�S���ʔܾ����M�!"������rO\o�)����g�=�c����PP�N�$mf*�������T�R)+�acW�:���2QB�N
!�5B��K,%��ND��;���"uۻ�>�E��"���6�f����:�@��NY_#z�w��MМs��0�*�U�U��0��"�t2G�=V��8r9�����Վ8��u�����^O�q[��B'�������Z����Ҷ����
��|�?��4c�_�;qFk��|Fw�sN<q�>�Y���⧠]���n5�DE��%��l	��s��z��hY�J� �N,6�}ϐ>�'��M����	�jG�8��i�׉:�Jkض,�;�/��s���L��D�%���p"�9�(n�*�漈LL ����"�Խm��^��}���h�%�]]#�L5.���=H���*|j��X��zW/���Hٻ+�Q0*��w��Y��}�	
�9m�a{�u	r�b= �{s��Fq���!���{�:�� D�g[��Wo���bXԭk�4�f����]k��5(TA��u�qj���h��z$���x �2���h�	Ǩf�X�;���^�Xޚ��iN��um���U�����U�z����N��>�҇�ae�W��ֹۻ�l[J?HsN��C�&�u�"�|�bC�״9hVe��	�����{�|p�|�T�a��8�*Z$�vL$Z�ω�\9Ԩ��<	&�`l.��#Y_��ޔ���D�Gt��/V&n2�O��\�l��/]��9kk�Z�"SP���;i.�媅�:3|��ȺX������Cӊ���$2����<����f ��yn�]R��#GM���2L=����3�\��:%�+�C��X��	�M��;,G�{��lc�<��ކ�/v8�����L������D|�HJ0j&�7�'ں����a���Z���Z6#0k*��]�����m��05xU!��a�~:��%��c�۴��2X�j����W�����7YD-ҷ�/�����,쁉�����F��V��Q �u��~��Yz�	ӇT��%|2&vROh����K(β$������C!1��G�) <EK8-s�gޘg�>;w�S򬲾�gi���k���I9�^#-���qo������ƈE��_ޥ�N��L�X�G�ٺ�*,��=�*���6�]��E�Ƥ5XN�f��L����<Ri�� O֚�>@U�P����`đ'�Z�[���5"2��l-�cQ�0���`����VE^JdI;���B2��6�apg���z}L��!�p�r#[�vh[���?�E�T"$Y�4�����g�� .�S\�n������Ш����[h1i崖c�CY���7\0��g��&�MX��(�>CV0S�*���SW_�F9rO>�d�ؕ�Cb[��hd�W�Nk��o����X�{=�kr�(�=6��z��(
�$�_G��i��P�TRD뾮$�oz��`v[�I��"�e��V������cLZJ"@�@=�(��@�����b�Tk��g����VQ��|�y�6�m�����Ώd��������h</6,�=xr Jo�U�-Qd�x㶿������7�f�3&�"��So�Qs[Os�>}c� Tق1�h�e�Mzj�9�3��ZB��i�$_�q�X!2�aތ���l1䋥�������P�
�7�^P�
�$`c�)Ɔ�͵S��c�Lb�F�q�� ��8�l��w~��ܳ��Dx���#][�?��3a��&�
����p��6��"�Xa�
\���ľ\o�1y������=�H��¬��S���M7 �c��ңe+��ޠ������ �ZmO��Rm�Ķ+�q���KE�,L^�ǚ��<'�OW�����1#Ԉ�~S
�F^�C:
!Z���q�� �t�R?0ۨ���:KU# �Z0��[�4=U���G`�#��Y#���m�����-0���j��6�_����WM䎮��pl���R��F3�z�T,y&���	������>j;�<]�b$��U�C<�%Q��ӘP��^rCUJ7߶t7�K�5��`@1�TR�e�n-C���l��\vFnR|�z��������-��4Gi��b`��m���E�.}&<����㷺OH�܀w�� �7�y�8��X�f��Z#zq��S!�yq�a��B�(x�쯶K
&FA��M���TS7������8��M�S7P�PJ��^�|��/RK�_���v�G���N�W�$/R�ו��/{h�;(�Z��5�r��r�r�l�;�9�¾�M�ט-�9�4�,�h����ԔL��W��/��	s}�����-,��.���w�镀�QtCbt�!UL�<�? �a�����~_�ވ��"�oG)���M�`	��Q�Q3�b�EԆ	�o�4]��]�6�p�/F�΄�VP�~�c`+��r2����h=���Q����\�����N_Z��GOavk��);���mCȧ
��\=��V�&����US������T��脾�O�6mjt�'��7>;@�����>�I����՗E86�	�Ӿw?3*��������4��'����2��_�܅��H�{��C�f��0I�Hsb`�mf(�8w�N�W�fs��a.+mh>.�o��,B�(*%i��װ�,�\喼�52�.�T�p4����v���e�!��tFo�C���q�<��_�犯"��Wՠ}�Ne�2F`N|��f���R���CB��0���15Lt���9ug}��T�P4.L�T���4��ꫛWVy�!�S������dz�aZ���w�oN�������/nX�>��c@��C��L8 �F�1��]�����&0�[�&ʫ�N���JUl��z�UO͵Z�;��1���
 #��bSL�k��ڴ�4r��Q秭_Ŭˋ)�붊4��S�{^]��Nx�2�D�\g���e�QL����.ۇa��;8�����"l#6�5UL������s��,�Zg�K���!0�SI�GS��qJrS�5��
�&���&U��G4`d�(��X ��TA�ٵ�r��&up�V������<����8�/[uZ�7]��y/��	�;e�8" -d&��l8�Ulm���s`�A��ĵ���a�@���H#{��js��j�tn���CU�-^��$�ز���������O�N�SN6�Ags�/�j�%��9d\�9�����)S���R9Ξsj3��$���Ay�x�諏��E��:�����\2,򠓎�ă�ֳ_�-<�۷v�ٗ�e���<2��wk��	0{��Q<.Uy��BQ)v1�a�$�Y��	~��^dV�Pf�7�w�}��-+>�h~f[R�����Vv��R��8�8�L��p�:�ag91���cS^�ļ�$X��-z#5.�ɂqr�
�,��&���ރ4R��+�C.*�5�)@N�����u��'(-#���d�ʒO��%�&�5��8�T��䒫��8�T%!4)S4�(���*�Y���!�z�Yd����\��ɐ[u���n�9*[vg4e�����*����t>��3�+5����������רw�-{_��9�G2^7[-|!��gaڋ�b�Cr*&Q5����=�p�H�4b��z+k��f���㱺�6%0�PNu����B� �ׅڟĂ|�%��^��Ԫ�`pkG����1_Z�/L�Z1
6�V37j��X��H��I��ť��XuV�rIo�8b���Q�Cӹ�k�jm<��B���9����,�ZP����;4Sݱ5^��F�+f^�J� �9���.�+������:-�V�b!�|o���*A"yAη��A��W��tw�!8z�u��e�8 ����!� $��ʁ�QS38����X8Z|%�]�(��y$#u�q��i={|�`�U��0t�LK�_JGAe�U#��Ĉ�_�hi��kOm�&�����&�]0EB+h�&���V~�!Fj��,	��oͿ�wD|���S���mxk����G�BӴ���ME�j����^�S�����rO{Y:.�50D��@����"���F O;`˱v��ٓY^�n��\p2*K5=.���|{��9����&Q���RXb�e���]�L2f�l�rS3՟�SS걪6.�wM����ڙN8{�� �a�?�� 3�Y�����Ɇ/I�	�����=�l4�x�~p�M��[��w��+d�%r����_��Q�[N�acfl�����'�roS�7�԰����rX]x�%�U�*�kv���m,�ۉ��[|���Z��?&0)}���,�-?9[�.���� �*�cHx�a�DE-,��h��F��9����Vr�DAq֛{����n���S�=h��d3����/� X4�h�\��]i�E�m��#d���j�RJ�.ݜ&H�W�Ɨ/%�>�5w%�t�ƚDC�нQaY�_<����ʲ��DE�_���>�u䁝iA9�4�J�I�5k�%D�o���ӌp��������A�Ą��~�t:aԛ�Sh�h��[^����Z��\�,��SO�/ J���R�'��8 	�nr���T�'7	�,�#��OcZ�9��](�x��gSO�-���v�B��.���J�h:`��o��e�s��;��˦!�k��K��2��m/�{8ύ���{�aQ��+�'�g�$�c�.�jz����Sb!���e(��Ƽ�b�-�4��rK�f����Z:��i_�!P�M�P��6wV�a����	��8���4��A�b:;�E.��Ǧ��h��]�G�#&)2�F;�%
��R:3��@�dqe�G$�lCu36�Ϭv~�9�p� (��-�IΙQ��q�#��F�pL��?ACasiӬ��-|�N�b��x3+��|偃a��ۇ�|��ᓘ��[3ӓ�[���y'! �&�)>(r�#�1�Ķ��E}��#a�Е+4��T
oĠP�rcn�H����v~L�&'\��ۊQc����0iWt��B��rLS@�{���2�*��B��D����~��kB��/⸲c5��t����#�����/c��*!x��RTh1�����-��Y�h^F������v���.t"6��ä:����SR8A�MQ3'iK��s	��'\En������}�V�
V��#���%Wr ��$%b�d>�����#�~*�}���Yţ7��WgZ�o�}�żHd*`}����#�gD9���-���@'�{6�i1<V���U@7�^�`l��S ��+
�ǘ�qPDG�0,]�}U���6���^��!��(yX��낀5���	���y�7 �����s�fJ70�ǉ��|/X�,��X��h�x�4=&0Qs|1���l@���y�㲒s��e�5�ʽj��b��`#�����0���1�.�*�&,\ǖX�Hj��(ζ� -�P}84۷�,[�Q1�#԰5w�ȗ~��C�1=�Q͟�b�F:�^�)1Υ��v�������N��V�������նV9�����<x���&��s�4Zd+	��t-��
遚��,=˫c��m����V����i:�0�V�(B�2CL�� �>� ���t�];D�U0�!�>�p�������@���*���Ն��L��n��K(ql��B=������q<-Y�Ng�g*���$���M�� ����WYᎎ�s±�jɭS��r{p��[\������Ǌ:3@������y�:���:8�^����@��^^j.T���QN,g���g�`������b������?{�>�[|Q.}�g#v���7����@硆bwߎ00u�̮HEr[

@���e�m�+���� s�[��J��s�E��A��R�ո�r2�0f�W5��n�<���4kW��no��t"s$��h��Y��_2|׊iR���?�e~�S�?�Uh�9��jX3��:���Iz�� �d��H:���d T|����r{���G�F���P�����e�K� }:��;b��0X�rm��4$%����"*5�F����$���.8�O���>u0��"7i�oHZ���b�)�t���@���{sO5�
z5����%�R=�����f��>��d�Gk!�+:�)��"��j�q�·Ñ}�����_)8�\�g	"�B�9v#�0?nB�}���H�}M}�cGus�r�69�'�/���y�&r�g�?�`����/JX�,�g��9B�f���&<3T�� ���s�^�rM�h����Dr��$ ��r���$}�%�]Nq�;���J�\C��'�ũВx��V'�A}��1\����e�OG�`|���v��Z���306Y|���`&k��֕�)���)��g�(�N�5":0�ӡ��'/���'���M��8%�!|)���L�L6����ѥ>$!w:��pj$;E\�(!ib_�y�?0�Ԋ�T�
ie�!s��z��ƅDt�ٴ�Ht��GtH2r6C.A���Ã՞�*�E3k�mG,����H���l��/Y4R���1��vK�!V��7��2N�2ϾAVl���c�b�9^�:�S�x�L���7�l�`�[O�N���-秇y��{��<<Ϡ�
ݳ� �Et:r@Jm�h���G�+�t���4���;>�<N44Y�p����-��vĈ�u�ݍu^�!��) g�OЮ��C[k�jxۺ}�d�(�0��#�+X`�jq��@b�GD�[4�ߙ���O��`��K���-T>HQXlxV65EB    fa00    2920}�]�����	w5������B���U��;�����i���,MIA�6X�u����%��[;̀l��si�\��Y�y��1��[w>��r�Di_��&N�t�$@�>'�^�'���q���.���8���0?�����b�j��Gۍr�.�6�ތ� ��oZ�]�7�Xvny���3֝����(�IgA��5�.�|F����w��i��B�š$?*�`!�ﺹI�m����F���ΘZD^G�4�}�2:����������z�ģQM,��լ�d��b��|�ߪē�#)����H�>�xk����	kQBg���O�Ӱ����%����c
�,��(�s&��
	Dr�dv����X���������[W�p�ӻt�`=U�O{�UG-�ZRi��/����]P�)7%����#}��Ot�$��]�/�D������}EN�E7=仅��_�@n6���H�{��x|����R�)Ih�+؜��:�Cl�2�u��dݙgs m��L΄(�K����$mK�M~p�N�$�_iy[��t�L�LX�0��D��ED���!uJ����Q��,-�O��	@W�Z���q�̃�g��h}a����<�}Kd��V-*!�&��7��=" H�I��v+��A��jNNm�̸pg��@�"Y�
�������2  ��)<�$0E�r�9���!nq������\$�g���9u�����孝>D��SXPN#&6��u	�a���ޫh�ę=��h;�����+�ʈ�{kJ������b�,ϙ���Y[%�粺 ��D�J"��@/0G�FăG�bU
 ��>�-�A\�ObË�D��Y�XM.�(�oP5��@#)�z�1��
"	��I�������&�UYj�BJ�ݙ��0���K�
�'��[=�N��-�Zu${%	�Mv:p��%S���z��X�a���z�j�� �g�,�[�H>�*��9~P���STp��$�ƣ�Zkt�E��։����/H�)
*G�ً��,t�n����H����p�K�$�Gh�f��#�FQpѡͺV�@Q���т����n%.q��[��\\L�JWzb1�Vޯ܂5���(&yZ�I�J�S����˂v�	1�̴���5k.��L����2��B��d��5�% ��O��/DE�؞�|4�&�z�#�Ζ/���%�E����ˉ���G�n���/C�x�u�@!���9K��?Ш�1p�nx)��.-�d&��� �Gf�Q�[)����D�wi)��U�&e�xuk�q��V	^9mE�����GfԷ��N�LiE��t�����ECn5$qo!u> �L�Q��Z}W�Y�o~��O��k��&���n�̑h\���W|ӂ��c��M��I��#Y�d�� cn���Rt���wuZY�ww�M���z�$q�A0����,�ƹa�|�>���׸�> ���w���8O����
���V�ۢ2D�V�Nc�n?��_�Z�'��G�Уl�Sqq����봤w�P�z&�{��k5XI+��\����e��O=|��=�lQ��P��K"ko.w���i���>5� pl R�&���4���햰�ӓG�
6m�Z�"\̑�}W�B4�R(����=B�:�������8�84��Jų�zm-��GY>:���b��\�Gm�QYz#�[h�rJ'�_ �au�$�|*K�m>������ѢBP��F�Fm���uXЇ#�ٚX?��p�)�G���?шp(} Ʋ��(�M�;U�zR��)ܐOV�^�"��6l��חަ����Բ�7�PM_�p�E��fg���=���y�@�X�o}���������d��xH��5��vZ�c A������#�vU]E����ʶz�7����O�|2 3[㋳�(NG����n�Ё��UhM���G�n]����QF�S��h�'� D�>��6���A�3t�M��0�$G��h�/3W�7�$6WC�s(�ǥx�#c�����4�%X.�V�-�\�K��8�*��|�������K	�<Y�����-y��`"�� #�!96!��Ї�)�/�ω^$��r+�E4�3����I������c�k�%���#>n��Q�x�۰���½�����@@	�֞[���#C�lٟ��x9�4)[|컏��z��	� f��I���ݴ�YW�FU�4>��L�����n	��[�~�k�c�@�϶�u���z�&�ӗ� �i���)$Gr����oЊz�"�����ƣ�1���J���a� �y�h7���yO�j���`;S]w���=�T!�j��#�n,)eP�B�5ٴe.F�z���p��q�����J��+�ܨ�Y�@%w|��|k�'��Ӷ�	���L�H�;�1ul_p�+5��&�[\ha�oJ$�\�]a�&	�.H�W��*b�h���zL��ЉJ���Ą�EUX*<�|9���O6+\_q��זnAʦ��IC�a�?"���h}qRD4�2W��	���`�n��N�	���v'�
,��(����^�qۗ(��_�����7��k�D�*�k������c��Z��Ȱ�_M����
�L�`�b;��R͈�>�1]GA���h<��m &��ל?�hx�y�TpNnE����N� l��ҏL��:>ۚQ~��J�:{@駻�(�f`�b/و��S,�ݒ�����Á��ewf�����&y�}�ƹ�8���4���DZ��B��d��fN�et����Y[�m���T=s�8���JW�N�Y�[~m���N�t�w�����G��n��*0ߡM�ѣ6'���Gl)M}Z�]*H����I���	<|�ӓ�Y)�CZM��u�9�v/�4d�.Pl�l��G"a�GY��a��Q��}׊��%_塺�	��TW��
��>���\Օ�*�.f�`��n#vjt)ܡ�6��d��AX�{
g��(]�Y0}���j���ϑ�{��y��l/�����.��ҀM���ǐ���6���J`@�,E����|�D>�;���:c�a��V;"ֈf輺-[5�� �"��ws�*
ْ7�nA��L�i��+�}pĜW�Jf��Q�-]��c9yk��D���UP�Mqo\�	=�8�D����]�4e&_�����n��G��ζ��-������O7�>��+�ĭ+�]ӄ�b�E����#��7}�%}yv���ړ�����y�G�J���#ԙ�Ɨ<���������
���W#�V���kvx��ve^�XĮ�jM�64��ůO���j�����6��ί���ˉmYq�Y
��QN�
4+��-�p�c)����%�-,���:���*��3����,h�����<:tM[��m���K��|��2��ȼ������3�)Qܯ�qR�C��h���L��°����)�����,>]���B�b 8�}��n�<��w���i��Wq�xM+��l�����c�]
kL��!l#�0&d�o!˧�����!	�}�Z��@��a8��jh0�W4eQ��SD�b�*�Ћ�2Z�5���(oC�	Wr��^c?�T.5�@�$��緘@�@|#5���d)=�	W������o�<G �:��O������5�����8���D�]ܤ]S��T2݃�KJ>��5"�%�;��8G��\�xѳ-���#�v����^��\��`fv\FH���WU�u�u4��7���M���(!�V���}0�l� ��:�7e['�19{n *rɒ=��(���}1�P��r�j�e�wRS��/�m��%%�GD�O1�٪#>��;L�z�!�Z9+="v�@�Vt�F,�M���|�'�7f��~��^����RY��4��1 �~�#<�A٣��g�N��CU'�=w���$��YGT%���u �@pd���s�B��y~��Sc�ы��p����W� 5�;J���0C�(C��Z̺q!]L��Hc�PY������� ;A���Q�FM9���b��ڀ�yb��~p�<�/_i��0�m1������.�V�5�^�8�RF�f��[7TmӚ�k��A��GgI[�f<���i[�'����z���-9ڀ#y̥�o���N�NܷS�('6��.�䞝� �p�MT�ԑ�b3SI:��"�9�]96D�1krg+��t�D���L���Y�)ZG�R�}W��Z�k �/�G�f
������ͫ{��)ys'�os���|�ݳ�.�/-X�i��:�oz��ٲ�a����țs�2� ���}�@��|p�y��d���Z|.[��/3��#�L8��ļ߃�ԯ�V�0�M	�=�wAeH&�'{zv���*�4����>�'���Zg�/���B�������V�]�ـ��-�w���H-k�Uh#��M�	�:�l�hK����&��vG�Fd���P�\S���g8�A�����P��Db�>y��N8���XXsC��)��P X-E"Z�&Q�
��>(>s,�&\C�l��)� p���&Ղ/��ض����&3x�bn�0?*u<}���c���1�J�hG���z�u]�=�E����R�pa넽�邙{��(��e�ݝyӮ)�i]L{�G��B:�(��ޯ�y����ġ�}����*Ҧ9Yq-~����c�O����w�y�j��`>��"���N����M��@:W�yj��x�Qr���V=�ZWi�Ѹr���=���M
�@_�'�Vk�'�\��ݛ�I��_Y9B��������_"p轼��F8�0xU1�t�>���HdR��&La��jzc/]�J�����vD	�l[!x��F�;2U� ���%��p�iwbE��'�
q�+�Ω#k�"��wi��9k�����h|�8HkǎJ;�F� )$�9~~D}=7_�E�:n{/U�6s$t����Ԍę�Vz��+Eb�(G�/�ӌ�<O�r\�岁W�Usi�=}�h�G]�&I�7P��9�QZ)��L��cr���y�M�#�
8#�{ĳ�-o}�������7eW���E�~���`3���і�Jw�*ԓ�`�$�נ�6����qͻ��A�(c���No0ԗd���>��*)W�2!��!c~�'�*�%G�6������Ҙ1#���0�(G?z.B	E7D�a[KĿ��)-���]�'0RƉdѿn��0�]�L�*
�  ����Ca�n@������?��ɴ�-)�G'-����><B�i��~dAfC}�Ǡ�sz�$��pU��n_ S�e��̽�Ν�J{�S�[�^,�K����;aU� i��|xn��1pK��L�]��Pආd��0(�ĕ�=��PZy����&�ts{��=]����킫�B�v�T��m�<�e`3�.�b>Q��F`PK�RP��m�c���1n[՟�� �����������+t%pP �G{�Y��$����롩g<}�X>��MP����l��I�H/�^�'��&���b�ѧz��>���m��pzi����b{WPb6� Mygs����oLh��R=y�h�h�� E�Y�if��p��sت�Y�g]��54�<6��ys�\�����7hbe(�b���V�FM��o���Tk��o�^16s��ƈU��aK��;$�z�����Hgߚ88�+�*�O�	z����N��[q4�O�o���K2�����U����r@�.\�8K6��W�E ڊ�AC��V��`}g�D��4 Y����:�|��P�9�;䉟k� 0w'��Ԅ�ƏWyG¥Q��u��*;E���e�����d=Wb����˂k~� C�ˣAԉ���x�����ô5����n����1C��##C�OHښ��m�qFg-�ɂa�z��y��ʘA)C����H�#���[�1j�M噱r���ɍ��t##�.�j���D��x�1�#�sk?Ӳ(Ev���[����N�"0&�U.b��F��-ցH�>L��4����p�[^�g�j��R����H���U��m�LPB	�.8��N yRo�yI��xQ�*P��v-�_nM�~JjQ�-��D�r/Uz�e26A�0d���ߜ���9���uj3^t�x�U���{��`�C/�c����U���Ѵl*v��(3y`���?��;�(d�;�4�m�� $~k���x�F.��}���!H9�$g���l�L�_�#�$'Np}F(�����գ��K�>�Z��(H��a�,d��1&nU[/�����p=Q��߀���
x���B�����#��%|��Ώo���*�CS�:d��I�
҆�8ԁ\���h7���r�Ȉs5��
�)�;c��9^:�e��7^X�m��#����s�ZK���v�HpEx���Ʉ�bCNÖ{'� �^�c��QV�>40	�B^Dc<�N� ?mO�1i��M���3�Ѱ��ˈ*��j�	� 9�[������8E�󨑼ZT�����-嗃����U쥰i��V��ԍ��B\B�{{����� �t\Q��f-*�(w����d�A��R)��r��H����{,�c��"��_Qn��D>�Ӳ��*���iKwc���ѷ�V��Lxp��x_���}{h `
�\
2F6�6]F���<�6�/�3�fz����U��/T�L`��g�'�שw���j����M	"׍*^l���"�7a�RM��C���/���w�A���<���X7�oV��5���h,�c�;��}tZL��MT���Yc�h��LaS4{���jG�:���lE�\z��l�u���(B��,��Y���w��Y��SƗ�m�f~Ϳ��d����0��k�D���܇�>I���p�H$e��6��]���|�R���i��w��h�����Wf{7���wA@XT��[x@F��+��ͧ��r��f$�wB�-9=���X��l&Xa�y&��(X��_�G�#�\��>ݐH���?�lX�γ�����J���P������Z��ʲ�*t?�T:A�~M��_����]���o�֮� �Kf+�'�ͦ�C�����69�2���C�����	?�0 �%~'ρA�Ƀ�����C�>��ɡ��P8Y�͊9��e����4��}u#��rO6�q/g�ݝ���K1<i�:R�r�^K���o�O��	����j��R�|+�C���e�8�=����k�p����m�Fh�y����6vH�&��Ab��ղ�	���"D�ҵ�ӭ�NU�,�q�F��c�$L2kS?j09h9�Y��Jf��F.�<��+8��;�]��o�W��H�bN�ag,Aё���v<lzYLPL,��6��&)�\���,&D��"���G�V6�9�
4ZQ��ҳ��4�Ӑ�� �k�?�Ƴ���T>S=��+rR�Z�="��L	628�%��ؐdUg���������G����*W��͗"��zE�l�־P�krY�K�� �������uG�!kf,JM�b�Oݻ�TOD���7�@#�>K�&k�nE�ob�R�,���EpGp���ϟp"r3s�τ(}��5��Ϳ��B�T�ӄ�E��d)�����y�\���H�7���!�\��;-�"�`W��Ө�H����?�2�<���rX��p�����ōM��p�i�'s���(�#^��k��d5�Sydh�ˡ^U�S!��'
��"ۅn�i5J���7~�)��ͫ��ӎ�8��f% :.�'q�d��	>�@2b�IY��RB��&4�͋����Jn�E��J��l�䍾7�М�?|�����xU��G��9�*Z��`�,8��"����щ�<N��GA�}C��ڂ��PǺ�H��;5�TbhL|#%rK���x��B�r�%c�����L�F�E<d[��ףQ���LE�����?�������s(xD}V"����tЭv�4M�T���T?�mԂ����gd_�:RQ�B*ȤcӍ!��]!�V�	'�Q�Թ�rbϗ��;��6-��M5W�������x#C�(��&{�s���2A�HJs�Z9�ƍ-���MīC��Ԅ��b�̊��*"-��;����9��M�nGv�$m4�!K0�Ԥ^���3�]w7��Ʈ������,��ėޞ_l�՝,s��[�{��УJ"����Bt-�ҕ���O)��E��0泧����?�w�]���G\��|&��E�������)��Q�����{�Y��Psf����i�N�<s�bMځ[�p�ѫ"�"��`	���L�p&���%iKOf�J1K�Q��З*WKy���`ta���3�ˌ�V���#l�Lo����Q��H9�d�7�K� ^8�ߖD �#��
S���$:���`QR{j�f�ݕ��^f�x�>��JϨi�r�OQ���M3��jJ!r������i��-��l�yGe�^Q�|�5@_i�E0_�}-�	���s~�vǈc�Ev�N{��*�!���e\x�_UBn/��`����x���$�P��M�ڊ��k`��-�G�{FPY����߻�nB��I�5�|*�����1!���퇟bJT��0�+jJ^�t:>�a������2�1>��BA`_47����ıݜ�cB�"��$�Ď���|7ה,OÓ�Y����>I2��v�����V���z����0j1��Vj�ϐ��pl�YI�<��������s�I�h�t���&k�lwAة��j�PJp}.��Y���~	��O�MLg,TH:Uk�[�&@;�̐��jr���V�U�Z�>H
\ 6�=yZe6���V���=� R���9nx]nc�I&�*�	�UhlV�znA�Zfc����4jB�`�s���3=��z�٘p�>�S��;\��a}������:e����U~���'#T�;M8�TJ�I��T���i��P=�d�>	�(l��Z���è&�K���?(DWW�$,���� $7#r~<���.J��W2�ġ	���>q�fI4�!?9Io�d��w�set�u���
��h�?Z�<�]#� Us�@�e
 11/�q����W��5��Rċ����9��6ⶍ��� P10I��t:"'8R�u;��3�G0 'Ÿ��6����X��ԁ�:��@ݡ���6`&pxL�����Ce�M1o�Y����R��>n5�}���D�1n{$:����L�8�LO=)E�CI�Z��M(�dW��[l���A���Cd����)��y_��ڠ�0�b:�:�6����Ƅ�Ć��.M�$��[�ji��K���Xd���s-���m����5�mп	9��Ա�BD�Q��P�^���0P�� ��\<�!ڻ��1)X�?�1XS��?���O��L<��(�w4�����el��*:���TY��h`���9(sq�z���}��$h�◤�@�L�ݪ}��df�j~Nj�Ȅ��b������a���FȠ�F���<ک��a_<���KҌ7;URH��:I������[�}�� Ѡ�j����*J�r1�݉)��¶��隀���Wp>���m��v��]����&M���(y�j&^�ˏ���^��v'�W2��ڔ�:M�߲�=s��eR[w��q��������ھ2eN7D7��sGx�`v���a�Ѩ<�񜫁7����џ�0i~:��ںǾ5z"X�̤���/���.������ �L�!^��~Ɖa���
@�t�eq.��Fe�FCi���+�~ o�9ultT�o+�} ����d.�%�#�Ox�Q�*S�?���3�9d6 ����2�� xM�V�Rد�
8���k�o͌��� ��E1�r'h0]ѰI���W�,�0>��X�3��ÔT>�� ��ق�b��)Ҧ��6Gz@���K��\i^��au�<.���:e,.w�FΠ�B�:�TQ�zj�������Gu�:W�Z�
5��5츦��uJc/|��$�Q��b�[������ߛ[c0���b��4�a��K����x�yI�u�	��z1׈��c&'�J2E����k���*wV~��bBKMb/9NXl#������c`��_/����&К�3.�[�|q���5�W�%8ok!��c�U6�Ů���qo��	}���U���	����;y��cz61t7�~��&FR�'sF�i�qL��kV�8�6�Q��9k����v	�~Ʌ���j�<S1dK����˂����S�bjz�*؂cT�H舐39���$k�~�E������o9A�JyM��̉<�v/9�!�T�Za��$�]
�&�� e��g�'x���e�;j|��ZR�)��Z��^Q쇿O���5����8����	���y"�%(�<d�e��F�4��CXmg���")%��3\�[�'m����nyn|�7%�"d5g�Dq� jZӜ�=���~0�	�b�L<��[�ѿ�aXlxV65EB    3deb     cb0�OMY1��I�E���^h���$�y
X�Clx�1;�Ϸ3�?�Ȟ�h��(�q�r�!'P�:j��`��]����f�:p�OW�ƠWG�$��x�I ��eK��D�*/����]�j*5�s� ��m��Xh��:�&���}M*��B32�����u��!�eq#
F���_���1���˳�I-�J��0'�M��Yċ���iR���$��d��})�F���� ��X�ͦ���Od���{�!HW( ��]�2�{��0�(8���k����#u�S~����X+�w�~�	�s���|6�n������aʴ�~񣄉5Xa�/�m�"���{0`l:��Ny6/xH!�տ#�t��s�^"���O0�(�h�$)��[��,I����mO-���T-�w��e�\V����K���~�.p
��e6\G�!����1�?|�C�z�,
��W&5�#g\n�����J��b�}����R���|k�Ib
�y��G����Y4>4���f)���K�*�IhsYI�R,t̚�8)���4���:#�u�?r��$PN��/�������%�a�����P$
���^���Fܭ��; ��vo�F��˖U��fwx�����G~'܁���j��
|���� �J�P���V���)}��cEbx�sg��In^�n����APDz;��HwX�B~7
�v+�0X�]u���z]ѯ6�&3 �-}r��
�i3�F��$5b�g�0G^�
�K���#�x�:���`Lp�':<�0�+A� 5ѐq���C���%�.��>'��.��o˦����9ON��p�xV즒}�vl	��2Ͳe��x�͑~kMg<6��>9�� �ZNP�&X�h	���3t�	!A��T���ğ��s]����\�)}�Q')�@`���9��7�8@�Ý�ڋy 'l82����R�oH}�{���ܘ�|�/��J5x~n2��Ĕ׋�m����ׇ.b��b���H��:S��m�B	不������7kݨ�'�2�i�}H�9�~�J���c�3C75N��ߌ��RGY'�#9������4�e��QTϝ5u+�:��rp����Nۈ,� ���O�,����hK����1�?�7���#��=��ȋ9�T}�[��L��*��||����'�m�
c�ȑ�H�d��Q�.F�=l���dk�]�4�7p��r)�̬�b�`�|c4\$�aL��H1�^��?���~ެ��k��T�ѳ���7����#��6�br[> �}x�0�i��2��]b~uf��q�P�N����5�ë�l9���.A��;o��~�=@6�]�/(�W4��2
$�2V�%��ɚ�o�eN�Lh�
�tB��XCs����q̏h���FĄg�9�Y�N���5�m���w�%�lKW~�SpA��>��Vd�N�Kةv���ԸO�~H��z��>q���qx*n�@���7��x^F���}W���̬X���<mG�l��J�ϰ��͈���+�:��4s�J��p�Pv4� �~pi�L�w��'�q�}���R�lC��-)t���j�;D��h;}@�'ܢ�Ek����=�-�6fܛ��ڤ9����ک�_W�>�5=+I��a�T�j�a��R	���7����d�X�ٰ�30��+�]0,����Ob�.bm�� O�R7�q���`�*|�o�kDQ��x����6}HA9�n�)`��g��,s���CS  ��	_��v���K#�ّ�<���t�c�H�t O{`�^�_'�Soq��xܭX.�I��;��m�w`9�v�r	Ɔ ������X���lӍ�hʮ凲���f73��Y�P�˿��Y���E֢�qVea@M�Ǉ���Wkڊ^2��#Ap�	�C#4d���Þz�4��]CCh�+��L�>�N�-��嚨-s+n2t�.O0����6����:8�K�atؚ,�rv�lZ��ʛߚ�T�M%2�^�9���w��F�֦��Q��lb��q}�u�ͶF�q�B�ͪ���C��ˀc�F�l�и���%���`%�S�T�yW��|W��:Q�h��:,�;���1 ,�c0�/:,�纑��P=R�B�O/��r�DC ȮF�9�@��I��0�7�Ёq�!1�Z��*�Js�w�����'���Vړ"��z\{�2*	_E�7l�e�`޲*G?�]�v��v��/����#��y��U�y�و[��X�q��<�b͔8"H�z��3���|����26;'�[�b����y��vB�4^:YWJ?nk��r��n�JL��`"��!�UŻ����ƻ'��؆@d/L��7��/�E�}�.c��7y���x��J��~@��B冕�H.�6��b�IS��Y���E�ѓ[�T�1���ۛ�Z�T�~H�����H_�o|�H�w4��V&�8��%�}�O|�O�a�p}���b�����~�|+��pb5�tTJV?��
��3�^�(�"����,c"�H�N���/p�=�L��ÿ�H4�9�r�KFu�d-��T�8ވ�T��:��D2��*�Z_*0�;�E� ��������-�|����M�Ek^$Cq�LK����,����[����1_EtTi�3Y����wӉ��� �|9�_fPI���:BQj���ܱ$1�#X V]�igwx���i٭o፨��A1�+��]^�/pd��ه�i�}���(GD%��Ơ�?y��wv2x&�q�TwVrS�&zYl_!m��b��r��D�sک��:���"���?�Axf�w��n�#�\�_J�A��t�KƜ4�V��P���(�T��)Pr�s�t!����Eh���^�i�dU�ڌ�!��Z��qDʳ^���}���Y�>�8fZBЎ��@?E_��Qb�l�B�Q����u1j7���̌��ќ[�(�hd�,���`�������pAڮ�s��^�O���I)�Tr�#��c%5g���GT_��2&'(\�,F� u���]�آPDo8�����;̶ۏKq��U�aIY*S�ZܽU͍|W�wk���
G�_yl(���{� ��@����FJqG~��E+o�/-G #k�cS���w�@�FO�wҒڂr��J�F��F��h�� ���ɍ����aIq�?o��x�$F��N���[�R��$�.�Y
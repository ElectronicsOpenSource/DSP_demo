XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C��Գ�I������4��@�j�2=���j�LWJ%O��w��������o��r��b��d�P���N��~�>V%�b^�ц[<�c����rd����
F�g��I���K�ʅK!�A�QиE���ԁo�;2~�Hܭe�ee��7��#2w�-N[�.�₶>
�O˟�j�G��y���n�B��Ψ��ᖧy"ř�t@v����"R�×�][{�є8�o2��J�I��zg������'/��=����u��2�"w���o3Dk�	�Bh|�|�&B�*j�{'�"�\�md�u��U<�@�i^f@vѽ��C�9V�M\u�.�?��&�YD��(;���`�=:�q������Q��&Z��<�րMB�ƫe2j^-�q�"6~��Z�b�u��l�AA���c.���-Z�9����@����í��(_(^f��*u����!���~��pt�]U B�b�̢�?̑�{��KD�J�:���u�]ycЪ��[m����9���d��	@:�`�^�M�4�i5cĈКK�����#�`�V[!��e��qM���N�޺/5K�u�tn>�qUd>[�v�8�'�p�BA�]_a�|�y�k9��c(���Q�'L2�YW'L�8p�xӟ�kH@C�V�1� *x1�}!��9Ns��7���ƥn0���D��[!��7��l�wʀ���䭶悜�-0�I�
��Z�EDb/��pjS~� ~��)��1,3{�sD������s�ը;�iXlxVHYEB    17ee     730jf+� �8tR��KP;�M�7�ٮJ�M>_V_�K��H,��r�w��*)�����/(��D����T�i��y�sgV�W>�
)N�M�q�ej���xjƾ8�"�/��u�Eed�GDwq�F5�rk�x�T7�;2�6�?�pkႡ	��-�
>�e1�֟���_F����ܬ�"	B���@�I��|�%0n�Ҩ@�'D��'��Rc��zh�x؈%�E}�����丮��54Rw3�	p���]�{���prȯM5,=�BUR.��9+���P(�K�<A^v(�^��/��$��}����4�����`�9q�k��J"ߗ86\��]�z�KR�v��}�Ny ��5��2Mr��}���t�gYW�"&��=����
���t�9x���;bv�
��3�Ee���;�g�+���7R5��$�I�~�d�1l��<�eF���!9��7b�癏��z^��W��!�ݒ��>�\A�+l[F��ڸ����u����l�w�F�$��ea Sڏ|Q�?����D/}��.#1�E�N�A�)�->��*�l��2E�k�]���O�N-�R�
�1T��T��	:
��NvI{Ql�z��b�AGq���Fǧ+��Vu��R�a����l��!s�x�D���`o�X8��^�%-�;ɘ��g?��
��'�uh�����{��		�"�W��Z���pr�c����{ �����]N%�Ƃ+�nZ+���2�5ѕh���������녪|���7�I�o4A
�ʾ��,}�����U�i�2hf�[N��[��J��t���_�Ɋd�6^����ȴT��#ؖ��Α��{Z�+�!�G�U���+����\G�|\2NЋ�!Kh�����7�Ko&�@s����<��;�D�\��~���A�^f�S|ǣG��`r$����Q�MQ�8l��K�+��b�L��;�a
fE�����5A�#X�yi��w�zeY�}{��@w;�O�ė�9T7�-�Csikf�D����`�^S���0����W��`a�N�V���:z�tJ��^i��`H���c������#>��Q��)ҷbL 1����7��]�� 	�Sȫ�3��X,��"�Uf3r�_
gZ�D���O��vmE�\��Yԏ�pޓ�B�p<�D$˃�o؄ �O�-/'��qEՋ�X9"՝�c��H't&Y{��";��d�{�`�Џ����u��`To�5������#���OV�����Ę�����a�z� s�!�-T<u'���vI��D�_7g-M���3|A�S�1&�~%Nv`��2m�=҈�#�mt6���M��H3ՠ�
/�'�Y2x<���������C�������(	Fw���#jB\W)lTW���+�������/3y�b�����򺏺��bn�`��A&G���@i��{r�W���gLd*���؊8\T@ܦH�y��Ӣ>(/�H��.$9�u�����(y�݂���Y3TS��E���K[E|���*~�����Qʗ�Ώ�N���{��+o������q�y:��eA��X�S�)��X��8Y�Lb :��R3\��(����ʟ߂�*3�~�����&�L�MgN�'H��zQ��{�������T���=P�a�Wց�T���q�Y�{���oD�ٸ���c��L���ϠC�m[Y2��W�F�nc�@]�0 ޽�0��}�.���km1F���p����nP�f��afcRQ�bP@�c��^&r~\�@��E��nz� �K�fR�|)I���^�}���+`Z�	o�`e�C,�]��T�����ٺ�{'�r��]Ɲs�;�~�
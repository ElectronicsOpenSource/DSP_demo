XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������&}�	i�ʵ�W1j�[P �t��G�P�<>�'Y�t���+�.����f%�G�  ?gr�;���Ka:�������n��Q"�����y؇5�����cCI��#p_lz'�W^�%�̿�÷uit8��rζgz�->5N��f
~��,��@<sYyZA����Tso6�w��޹I��/��sZ�K�;��I|hഃ���Uv�k3��sj�]k���\j23{�3�
�I��2l!�]8f��1����P��J�Ŝ�}���Ɵ�{~x|�0w*��9p��2ḌC&��e͇qn3NQ���N�h��X��XP��T0')��PR+���67vB�C�a��=�%�P%>�Mc�1�#xE!�s����<;�$�l�U)7�!����P؇C�eP<z-j�4�;� ��Z��;�er�j&�y/2�ҡ������m>�s���wH�׸_�����[�嵇��s{D������9٘}���!�߈�;�Q����������ڟ������Q�����r2��a`�x���[=,3�V���o�}4
�`�ꯁ^�
��NJQ_P�MMO��~"���-�E��pr�>Ǚ:Wlb`��I ��V[i7EZr���`{��gj^�͆k�g�q+>b�ҋU�4،;}_D�1.`x�km	#*��4��F{P)%VϏ=�N�����\c:�b�L��q�`O4��μS�>�Xt�x���֐�6��Z]$�/����f��]$��(�X1���p��xXlxVHYEB     e37     6d0J]��f�	�a��'fڣ���;��2"?�j���SҶ��T�Ś�r��Nhrq��X*B-���V�aљ�������V�'�2���+iMx�QD^�\98O�ҋ�E�.8�>2�6K`�Sx���+\���7�Y��4���a������ڶҵ���yX$M˒�Rd�F:��p���u�9:�,uG���Lu���gQ'(�Y埡�q6�z�H����P^*:�MO�oPG�G���)"�d��!x�����6]�
�)�5��e]k�jS�$bW%5�6dׅh�[��b;Ar���(���e3'7��I�T�z{M�	UЭv��<��ي���̿���Mkis1��d�X0�nS.�l
���ĵ�Y��
0�*����$������<(Δ�$��u�ֆ�xV������'㮌�I�<����{����m��Ǩ-�	�4;J�1#��#����<vnt�j�{9I�Fż�r�eeڂ6�+W�U�.��d� F�
O�M����'��$���"]a3�	(�DP��r)K�<����,ד��.,H;�<C�X�uO<��}�(��~��GX��SfmA&���3X��!�9����`bx2ܝ�^\���i��ؾ]y��H��a/յ-:%��s\�D���z+\tZu^2;�ZM��a�=��S�|(\�D�ll��)1S�(C�s�����=���>h^���r��6��iD*�v Ӗ�mHa��1'Kn��*^@���UL<���A��p0�Ռ�	��z��+-@���d���=O3ݸ��0�۹�ʯf����\ƄҰ(�dȶ���/�$jkj��,��M�|���s��N�A�X;����(�~B/�3�ۙtW�{K'��KQ�j�PVe��\�'.k=�OQM��e�=yT)�?zR�c`��-�`��aj�tX2�6W]�<~��jzg^z�8: �X[�'��]&��y�a}�n�1�5a����ۧ��	�� ��S˃�C�pWI1}�:;���l¨�A6!4졲 ���n�Ԙ[��t�Bh���פ���y��4��[4:���0�qφBZ}�b�����Z){��;S��UAb�Qb4	n#ر\�WB)��5�$�t�Uo���0n�S䗖ȝ#	k%��v������I
G]~����#T-�J׵�[��GE#B�������w��@G �js4X�ߘ�X������)7�S4�]3JWl���YV�c�罈h3��My���&,Ƴ�'�?�@q�#](�m�Sr�)�h�ck���n�OQ�����X%�2�G��dJ@�P��F��7�����Ͱ�a�'�
�?܏&�	�h��+�l�V?x��F#/�-��z��T.Ĕ�Lݍ�����]��ʀ)�ک�T=����S�\��ya�����%Ʈ��5�6�e��ڒX��^��Z�k��}P�\���1�s�������'�|:�o�;#ӬIoLG�j�s@1v&܎�j��i��e�� /!b3,$���I�����hxU�C_��t�̩bIڭ؁lr+�:�&"�NI㌵���f�nN��N��<�kk��T4W7i{�HX$���@�Ǟy�5}
�������C{,1�!��^N?I-���}�dU�%^2�t=�}
��o��ήi������s�{����)��y4�x&��@�m��=5��fI�Ո>�j��$�=	-�jM�؜&s��s�b�i���$v!����#��=
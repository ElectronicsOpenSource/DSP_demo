XlxV65EB    404d     f50P�A6��l9�ny���a�|%~�����nm���V�I8H�d�٭����̑_�����H}):��W���D$0��J5�b��׼��>����I}ߚ��;��m�T�#%{��զ���L��38�
�����Ld�;h6�KR6)�k��B��{(�rJ�$�K���$t�p-�N�	�JK?|�Y�$Z���V���*�zr[*������u|3L�1k�AUg�B���%��~A��:�����VP��[맄k/o���d��M/�K�Li����x�.�b
� \͓D�2l��/KwZ��ė�}O�� TZ'zi�%h�ϷZ@��t|����1+�g��Mb�g !b�h��'�_�b�U"�#�/g@~^V�(�w �
��r���Зo�S���ʠ��	@�"u�0;��3��MH̘�#=�I��j����\"[S�I��U�4��� �oh=�L�mP!X�*X]�>��f��H�j�a�U���;�Ol<8C'��-���̏�l�6CQ.�M>��G�9)70�!խ6��H�Q[��	ׯ��;��7g#y+5~��-�,tY�aݚ�ع<�p�L�$�i�.���;�i��&;�J�$BY���w%�O�~5��V�q D_�4YCj�%��V�l~�S14�e��r��q�-���t�k�&k�Q��7�P�u��׍SkDY�)R��8@���9s�2â5����+]&�U����ͨ*��
c,���E�Л�#��Ryj{�ŋ�:��t37���t#
��dn��?��/��'�S�V-m��j���\92��;E:M�(KR]�"b�~���(��^��ؾ�[�nTЋ�t���:�vg`�b6�ۈ1���l��d�i-��]qU��~� \􉓁�q��]5
�.�G�'P��ap2�k�B�%�ᴁ�pl���B0,c3�z�lϓg��_���i�Hr�܋�w��UF��1� [���6%�����8�i`ܶ^��(�k����4k����>K7N�fn���:�5LZsn��=�W�S
�{����Đw2�~���4@��U4��o� EV�F*k.ň��s�q�
P%'��^<_	�:fp9l����-Dn_O*񹾢��Tw�.	A�h��mC.Y� ��� ��,����Yґ�^�J�d�H \y>e�9Ayn�HV?�t^���W%�a4�wXM~��$�S��<U�T~c
D�E6՜%��m8��\�s�5g�nUT�sQ�-��x��@�WJo���d���K
���4hʦh�<`̪G_�? a1Z�����閔�p���I��k�¤A��z,65T�������'qp[�}_ �Ч���,,���G��Uw���`�l�=��W�'�t�=��2ec�$Q�6�|Dv	��jn�G^8$�� ��D�"�[ۨ�EL٢q{��"/U%���A�@%�*ٮ����!��#"��_n����Z�#�,���}��b�mL>����B�eQ�>ДDpz�&k [()u���t�T��.^�bذ�`Dsk�� �	G�k�%X�W�q~JU�v�e�*V�K{o���i����`[��*�kt6���Ѓ�N���,�6a[�ȭΝȖ�;&�O���	hbt���!��J����U�>�'	9T��*�}�N*��<���<b
�EH��4���L������~ο��	�h.�r�h'�Oq��T�:���ݎo�֬u�TG�U	ʘ؏kg���͠l���)�������|u���$���rX"�65/:��Z{�s���e\�=o�A�-ȝ�b�@�+׫�mk��������z�I5�s޽򣶞����{P}���F��Ca�v�w���@_״�qu�%��w��<�q8�f���H���
Pv)<�R�%��FT&�~��0�Ӟ���G��)J �J���F�s��U��3rTvB7�MH�����4:S��e5XӀk�Ú�����+���ʺ��'�.j������_��(��%����i!��gUN_Ui]F]ѵX@�<��_J7U������z;���
��q�bt���I�b�4��f�͑7��P����
�wT����H�;�4�m(=�ay�bk���ʁ���G�Kw������|2����9���d�4�fE>[=��O%����1}�
'��3(�Ƚ_���(�*j�U�Ȅv(�~8\\�J�'��dp��N�
�	92�"^�4�]�OlrW������S���e�Qᚅ:G�̸H�HK'(k�1):M��ԃaM�0M���"kߞL��C�:�'��د@��%�T�۱Ά������pl�ʺ}X�� �cE�ߓf��!�(m��(����L�.�E���=��Y"Ŗ���qF��g3���#��e�u�Z��V`@~�i��p�TfXտ�/\ςUV�
��vR!��[*kk�; mdUpv�b7렮�͹V��y u�%.�� ��ǁ<�sԞ�y�@P(�a�?�c@����O�X�f��en\u�4\��h����IU��G���4!�3Lh
�wn�����k�g�8?�b�e�<�ZQç�0E�j0d\1�{�NTmD�Ui��)�H[礽 hJB��g�ߟ�a'�إ��[b�
�Բ"�F1P��"v���7{�@b-4�0dWu�g���n��5�� ϘS�����~ڱ�Ww�yݱFP��!B�O�Q,�!�qq�԰0:K����$�WsO~i�}�l��fUM��][Q.��7ʂj�*��o����im�7n�zÔ�k*>�}��f�3r�G�����	)�9����a]�s��uF;<3��r.8���2�ܴ�:!�겆/h��ED%ٕ�*��3���M�/q�v���m�f�+XY�Ss�n��r��'��b�K�q���h9�[x��U��뻺�(����D�Da��f����^����
1߮�r���NAz*7.i) ���1�:�y��猚D�خqF4�u�q��b�'�͐S�[I���+��)����<L�r���Mth'+�2�-�;���jN"��H�tU��Y�1Y�;���c�=}�H�^�Z��ZN��9�D7��������1J�5%��U����W���8�_�tc�1���ߪϠ�-��1+�.(7:�eIz�tk��S�l2ёP�n��̳�i����֤�Ȱ�і����1/�#"ٕ�P�Fӝ���x���5��~\��c�#����Ed�]���7z�v2��e��#�T�E��,�|σ����M�\�K�Mޗ��Vy�C�.K���6�"��pV�SDg�Uڃ�(u��dV�"�l �6%�$��f7,��)��@*�	L�L/![���z5�_r�� �g��[��8Î�[�ȳ]�h��)6(�_$��Y܎"Huv<�w������F#vNk��1T�6u)1)t�"�鄭��{�$���eQ�#y��rV�[Ë9�~���5�
��n��2���$�Z8��]�>qz%=o4�PM)|�H�1�1�%8��Z���ҿ���t-���jn�Y»y��WGtp�������g*��	�dw,���ضkK��~��ϗF*�Q�fKll����Г����r�D����/��2f��·U+ҲnK�z.��By��nSD��'ST��߄ . fh���Vq�6x(_@=ޚ�R�5���A}H��7ԓ;&
��l8�?��4��ð)�p��Q)3Є�����Q�J�*���s���u�#�����!ʯPN��:u�E�7�	j �Q�-D]��=�������rA�Fpj3E�I5�twԪ`��b�D�)u�h�:���
��S�W`�>�G-�'�=
alD,Ҏ�r��e�ʶ}�)�ڀ
XlxV65EB    fa00    2f70�����O(�v]����^��L�M]��\��dZ���NG�E�w�+�#)ߥ�+]������Ӣ}�����?��J���8����f��5J��0���&�^�'0l�#�앣#�<a�P��am�T���c�j�t����\F�_s!��X*p���� 1���w�M��}�1*<��&g`�����^ɤ�d�S��=�aO좛�9�9<0g����*�IE��5���@�?`�kTbz�B~�y�D(�����s��G�b�Ҍ-��k
o�ʤ���[�+M�%���&H�BN����/ݦw�O����e.�+�O�6�
O���NϟLŠ�Ĭ�Q���X�D̡ ��-�\=�@/�ե��1���C��y�cN�PN0o �X�o߽EVk���W�z����8,A6�_�U�n���:�c���'E�VZ9�:+��w���뭝�J� t�����$x��k���3S���/��DxtΥ�+2�_�-a�Wo!��Q�����"P�]L0Q����P:D�S��k
Wm��� �"�E��I�
^�+�ɫ�"�kY@Gc��ٷ'�L�&{^��ߐ-��Ӊ��uZXw䚵D�o\��?�wI�*�H:��˶�J�Da�l�\{�E���H�<9��d���C,Kh�e��Y��sq�ՍU��[t���10c��F�G LS>�s��5얧Z�~�; ��[��O�A��{�M�\f��@�O��2�z��)��JČo(
@6�Ԏd�D�0��O�6����9�36Z�:fc�#��q�n�Q�,�*�{���&���~5Zî1��+A�뼋���E\|�P,�X��:N�4M��F����Rz�����!Y�6H��j0�~�ھhӊG��r�;��YA7��3�[{��s�5u�V����&��N;l7���K����4���Q��7oE֕��w�@E�T�x�<`�;�pS(��r%+��x,q�M3�+�����z0]	E���=���pnSXS�ָJ�7H����St�{�{��p2%g|�+"H�f⩒�뛄rQ[�{P��C&@s�3{����a/��H���w
��$|R���|9�]A�j]P��/"��d�j�u%("�o�5J�W��k�B���pZ�G��7��c&��%��Gc�Wp/x7f�A׻2㣞S_����U)�^ d�7�����G�7�KE��p
e�Y2�O�-1�R,�zڊB�G`Q�������P�$pYCp&s�g�z�z&^�uwh��#L)��`d�/w���4?E�TO��!�$�,�+�4�L�9Uo�XS7U���$4�:iE��d����_-��o-1��o#�J��V�����x �� ���d߱Uk:qA��D!��t����xD���ɔIo�4�(5b��`�arE/��Ɏ&)�����,!4F�z#��[���H�!�IF��0�}�rH�0��2�������f��(v�]�b���y^�v(�-q��3Z�����t�5RW��%;��٪%wB�F)g}�,��ܤ�n�� �KN��x�,���݌�#���7
��ƆL�d=D~��6���:j.��ȡ�%�`��)e��)WBb��\k�7Q/��)�h�����u����a�\_!]D!� ;���&�oWH�[�	6W��W�P��R��\�\x���4���ǉυ��ր�~	B���j��E��J���߻��8������	rD1��2yKE�4u�+~R3_2�?+����؛�gӔ�l^�8.l���{���U��\)g�3/��5/Ha���y�l�OoCPn��[�,O-���C�N��0Zt��	9x�H"Z�|k&~p8ל����J�D�~e����)�Д`��v��_���2cz�9���#H���gb�.*߼�^�+$g=��|S�r? �]�ο��k�}�ꕫ����+��$(�&w$+u��a	Ѷ��M��۲����E�ub���	2����8aP�ݘ�?SN1�/h�������m��Ԯ0y8L�(H`w"`�qxl;4�9�J4�>'�'*L�H��lk�5$CF
ݾ��äRO7�����RsU��,��P��۬�X��K:�z���D�T-Ma]�X��j����>S���(�Wݵ 7g,Wd��~^����^��	�n�������o;z+A\̀$(G������W'qk���#�R[aɍ�v�|˪̕�.��quȘ�{�*�T+��/X��C��p(��u��V��#���������Y�ݩe��U|NF����s��F;�:�O��w�<K�΃⎓�M�}�b��4�!�/?�`bNz����g�o�_�%�{e�$i;�Q�.Qk��ZIp��M"[Gz���)��5����3$n-mT�t:�l١Ԃ�b�O��ے��:��p��{s��b^��h361�X
������(�B����<��V��c�pܯ���/��b
���%b��rT��i��Q8��kvn�Y%:�3���r!7jy�$5�%���Ca~�h�[,�EX/?�s
�N&�y)	�ۮ�6���۷�Kb{{�-g���Tf�����+]��g���aI���QyY#-ba7@�XҔ�P�pKcO��i*��r�`��=��C��	*�G0����(���so�5Z�+���Y0���"t��G�lJ�l��e@%u̩/;3��p'2:n%׆N��&��A%�R�E]�C�\�R�?C�z	�=��ütG@��y�����o�>�lq/��n ᓜ�����)ɯ HB��K�՝�+��<W�`���kA�^�L��6a����z��13�ƶ��Z)���3g�o�I�Qa�0Io�";���SK���c�P��T+�$ek'5�t��h���_�",���s�:.�B��-��l�5	.2Dbn�0�n���))�B�j�W�+ո�{��H�����q<]��������]KD�:�\����ʖ֞�;z�.��h��"F �4�H���T���\��<��AZ鋡�9�G�/[A"�jx;�� @j��CA��In����kX�g��ި���h�}�SL'��D?���p�[��y�dne�5󩻋�Fq���T:Jnk���+��N	.o�Y��s(!Y�������G��BNi��9�_Bd�I��� �P@�0%s�����m݋@��wJ�g�x'�a�#��/K��5D%?M!'��d*X��w���j�]+)=���L�ͩ�,'��	�'Ɣhof��h�h�m(��Xό*��8Y��פ'TT��lD�i�e�6�þ�A�i_�U`�,s	]��U�J� ���:��@�X���NHgf_pa%_�% ��������~��*��UJ�������NQ���:2���j�"�ua�nɜl&h��O��1	V�����:[���L�*$�ɗw'��40j�_�#��#��oC<��A:�WY�?i`����%?1�/y��"?p�
�Xөe�R��^v���ia� �}�y*(FYm̍�-��s��^ͱE�p8�x���U��;���_��y'�/��C?��t�zZ�PlQ�����F�c��kǖ[ڙ|N��1�(��dڅ�]���`ѷ4V�|Yc6��X��.�gޕj��I"�
��z%��\��	�yg�� �cM�066��~/��N�xwt"��,x{���5���麗��o�Р.Ԟ*V�؃��/�ij>�,�Rk~6��/��Ob��z���h���K�eQ���1�r����ǿT1В#I�H���Ԉ_i[����0l.[kE�-��.
܃[�"'�p
����"ϛc��O�qX
l�� �l��������==���BǹO_�,�⾽f'h[��y����1?�hCn{�E��v�B�$�"�a%=O�Ɛ�TT3~-�+Yӈƭ�����@���.�F�XU�=��.�ܯ�؍�?�|UBn�y��35��
��+1�Ο��8~�{^	�����PD�? �_ĺ�xzK��׽��&���x�YwP&2J���( h
VŐ~x[l�M=޽���9�x"
(��hO��m������%�h�)Uc��@c*һ�]�&=�f;NAq-K�&������^����	K�q�i�r�/�����`��ܮ��E(�uq���v����h�&.����h��i'�AXէ�{�bT����������fǿ3ٌ�<	�6�5 2P�#.���#r�=��"��#N1�I��w�ԭ/�13���-�("�,�#��Z�(Aetz���IZI�y� "�x�\�f�y4�<�3� q}zh�����C���7Z;�>�����p���i����֎���F�q�^ٴ
O�V:�$�ѥ�Rx
¤�D�8%�TbO�{wI�ZP��f�Yg;�d�XЌ7����N4�1��
#�ۋ��ơ�%.�ǥ5'�W��O�i�)t՝R��.�8��x�QZ����Z����m�!5����.���ƶ����� C�={��C������ܫUJ�w��E,!;�Et~Ђw��1qˑ�,|6��
��x�n����W7V�q`��
��������s��oų�l����J"�N\�i8�%^��I�D&$��>����C���c��Z�)� ���ZN�]3o���c9Y`g�1$�}�gZc���l���i��D�K)����K���x�K��u�Zy�'������˻'ͨI]L����V�vm�B�ԛ�=U5 iE���G}������%���H�W�g�˦�=({�L&��ǖ�� ��X<<e;PF���x�j�/ve�W�����*9�H��0j�=%����t��Ã* 5��腰~�[�|m݁��`϶�;�"�yl�y�� �a݈ )�AD����ln��� ��p3�oOI����Y�eI�Ƶs�½�>N���%��s��£�h������e���l3�(�B𘞛0��	�5_�����
��H���`R��NYε��p�c9�����hz�M1Y�£@(v�#$��9�L��jv/b��Fr�?a���d��<���7?]_guл�3I�YV䦝i�z	���ٿ�6�h�>�):Fb�C0s�NSU��t7fz̯��9��8/>ex�6�t{؂�N��0� i\0����2���,����L���-\�ًPv����}�l��ذ���p�̓�݌Ԍϻ.g��˦�*EF䎻�1vm�q��A�f:<�ӓ������GAy���H��A8+B�~0��
��p�Bʴ.0��"b�4�Ԍ؆���z��[5'�﫵)�ь�ٸΌ�t�	C>�T�I]�A�8�f�����u=�&H�UW���_�Ž$J�s�Z��rh�b!M9�.p�^ȍ�*u.�~� 6���ŕ�&x��9��C\W�ɺ���D��zNܟJil�-f~��E0�o�����-���( Y�׊�{�C)&���.�HH�ȶX��0��%sf���`t�{�
a9���<����� 	U����`"S$H���r�]q�ۊ<���Z�R�S�	�𔤺4."�;�	������|��].2�����&��W=��f�Z�x�k[E�'{i���#K@Iy�F��J�ĠMen#yh�,?�ud�.��v���VxE*V0D÷������#�t'zgc�D_�ȍwa]��C;�Ƭ���j6I,������m'�"B L�<�K,!�!����&��2 ��;XJ8~������w��3B<OI_����5mn�$���l���T<�R���2W��2$B$X(3��l�&��Z1G�ռu`�/
Y�K0��� 0$m���Q��m����n{["��f9LR���4�|�XOb�Df<9�UU��s���k&�Z�.�q-J۲֦�D��*�&X�,)~,�i�\A�e�;Q+���/b6� �q% wq��C�=��~�tͥ�����{��_�\W}�.ݽ@��+$�1��AQQ�P���xj�[|r�&w�߳ꌄvl�Y�ϭ���U\�?��� sы�̈́�����l�F��,�|U(S�,����椃�Ɯr����\� `>[���jY`pd*�Î�����mȏ�?+��,W�SR�4�,5[i�%�Cx������L�"���M)���>xA.��R#��{Qb�4�ȹ�h#���\L���K�@� [{C�UL�cA���F�N���M|��Jv�#�
�$�" ��HA�Q4#��=��f�f�W�[��*�6,�;eO�ߝK�?��zޘ����N�n%#��Q��Z�ʡ�"-k�	&y��8P\Pj&�+R�O�B��SN��j�U)a �.
�k̿��^6�����`�t��i�p z�JrW)	s��Ӑ3T��ڼ��oH�"��b>��	�x)�)����_`�V�x�!���x�O�U�Ģ2�S]���훗D���u�TP�_��ep��ze���?��;��#jv�N3F�wv��V+=R�5����
/֤Qc�C2�Z�N��&�-ʊ�����PgPHt'�}�$ "iH�Vy�gͼߒ�-7�����@&+�2��(r^v�v�����U�&���x(���,�h�����hD9i��w�Ĳ{��q�����ʩ��Y�����Y'���p�ɗ���v{t�:�3X��YtqZ��)v���=�5��0�RMF�V�y)eg�ioT�#A���m��	GH*�� o�����}_fDF�0�@cZ�f�aXe>��hp>�@`-K��`�r�x5���qt������f�,)��� ]H4�:�8���;����������n�(:t���c6��&��,O,WiĸBR+���գS��^!?�4�Rnz5Λ��Y��r����?�;����|{|��lPr)<�V>�״�&33b���O��lG�P�:�D1�e�
�#�ŝw�A�m��"�ݝ��Fr��=c�\.^��L^2�e���#��A�/�wH�
�F^��W�� ���+�5��C�UG4���g�t�b�W�3���g%����{w|���7�ʴ��z�LfJ�@Dm_ZǳR��5F���	7�G��㘊�pp�ZF��(i߮6��9�ySG��7�+���83��2H��%n��a��+!��`؂og�vd5�W]b=���!0����3���=ѹ���HC=o�rp�# ��&K��'BȴJ�� I&���5@�ʜ_�zK����^9`�����q��ʎ�ꏧ�IҜ-A�7pFŃl�8��~�H6�
���H�=�xO�KI���t���@`����Ai��Ж�aI���j�i����%�x3�Y���0��G"[)�z��{�g�5�(�1��C@�+T�u	��q��;��O���i�!$����7@�t�������<�(��Oj�G�οj4��M�H%@�J^է���&]��G�z[�s	�q�����	���YA�G1B+Y�m��ݡ⌽E��_�kZ��	�Pn;�cb���CXty:j�ǝ�u�����ʕ�(��85D��'mo�����ˋ��F� 1�p)㜢��8;���<+Y�ytVQ:�g��˝i��A�^k��]����y���9�H��tB�-3@����`��4�UIȺ�5σQ�a���J���� <��"|��J�T�̬�х����
� B��d��a�1(�ܨ%��&��X��� eYi�\���JNV'r��W$��o��=�n�νC�	V�;iD���S�+�g3����Ux)�9'�u?�ނ	8�Dr�i�,�`m^&^��S{�!��E;)� hdfD�O	�5�2Yܓ���g}��()���;g?��[S��@Z�	��o�n�䠤sLU6PK\�����nu�My0��fZy�u7���,�s4����K�2nk�E"	a�J` TOm�+�d7�6������D�m<K��:<�s�e֫ۢ�ő����r��_�ڦ~5���]���f��-����`���dmFo���_����\�G�1���^=F��Snw���|x�LI���C^7$�tjB��0�_�>����ݠ.zi�+�2�Pu�#q�!t�Y
Ȭb�_��q�k�~֭d��F`�|),):̲��胕���Q�d��<�jL�<XM�`��lY��9<��N@qϢ���A�k�&���Gz���N9�H$�ʹmMn�%��[�/=���xl�4lZ5U���������>4T��!<b	�;z�.>�~�+�Q���y����;0C��q��Scgmað(w\�r�*���@kp \:��-еi$-��{���2U
	�t�8p�2��gX��H��O�	J� ��y�{Q�n@x۴����w���{�HR�cdkU��;�y���'_��xG��>��.�EC�+»Gr��]ܦ��tme&M������id�\�8�u%cw�m*��;1��hl��S[Y{�W�3��i�L�3��^7O���T��i�S%Q�ȶ|^��X̔�s�4����
��3Ӷ#��F���C.�Iu��)����RxD�e;O��@�P�{Dh8	*k��R�I���i�;�̧ah��B$���b��r��)lU s��A	���V/�b�PQE��xs�<k7b��V��4WD�!𷎗t�v��Bw�uO(�҃4.���p=�|4�u��o��� ,��s4��C����a-؀�2՝�Dd&��S�q���.Ӛ��+�	 :��c毥a�ی
�F9*��&��f��/�6�"
�߿�I*Ro����3���A���?�e��⃁�&3/���L٥�4�7���}��jt}��Y��Ia��5�gdq'S�"f�.���	hc"�����S�4�*Z������g���O���g�ǣm,��ŏ���j����	�CLBI��~���R�g	�硁u7�
|��^�w�d/G�z|��%F��DZ�@���a뉈����7��+�M����5Uս!�f��|�1��[�[�}U����̍Ѱ�)�쳈d�#.���= v��e`.�a�-�f�dI���R��Vj�Ǿ�<P�����7��c�`c���ܹ XF/h�\�N��GK#�� ���-�����ۆB�\¹����n;9M";�&1�D��E!�]�*���w��~��f�-ez#u=xzݎ� �ٖ?��� R�;:E�%g�a�;D|�>�'�.oaij�3?�o��q��� M����,v�$�/'ԔD!�J�!��>�
k��WA���a�̽ϜpS�0}|&�)�f�]���a��@�s�1�'���2���ޅ�G%]/��eb����8QΌ�L�>f+��t}�-7Fa���V����T�����*�EL�s �������"�W�38��bX�8����'��ꁜY�e�/T�1���y�����NZ�&$�t:,Ҽ��f3W<�	@5Ҝ�aCjꉕ5���E���R ���,�w�<�x�I��w9>.9#t������a�o�كlK|�C�sʦ`�����=�Ʒ(��Q�� [�bյ�a[����0!��ư�6N�ˉ��ǅ��c�ym�hc���+�WF�!��z��׻���˻������������۪��Izۓ��mv���X�CC_=��"�5��,����CC4h��?����4����J]��]b�H�fy��Q;��&�j3�9�[���A"�n�>J�(�T5t����P�?� ��ޗn�┷ڙ����4��p�f�eY�ƻ�Þ�+�1*�r�<j�@�gImNf-]� P"c3z��7������st3c���؎�~?�9��:Ki�V
^F���p��9�'�'M	BoeeT0� ��N��I����+��
l�+���>�kqܱ	�R�o�?�cfNrm4]�o����9�!��j�+�0I��S����&c5O�U�tKn|�w���c��寿�$�Fx�*{�L� H=�b�c>#���O웉���K\���u
uQSC����(?����;�D�����-�D#�'+�
3�/B�q�_��o�o�4Ip�IX�|~�	#�G�����a�����8�M�u���H[9������$@@
i�毧�0`ժ/��3C��?R�]�!)뫖�%��ݸ��Q�gD��k�v��
���Mf�K����]qN��vQĞ���Nq�i��1�e�f�A�nk�`v���m$l��q�x�p1ɇ[�w�F�dP�|����f�޺(�*�:��$$x������ׯ�%�h��L�C��;�|��^�4yPt��E]Ը+�Pjg���H���vs�*�?�L}n]\dUg�,？u=B<ε�#��	v�I�!�DY"	�qܣ�:�YH�g��nt.\��z���i�����rjk���jnZ�����#�� �?'��/ #]X��	>��|�����=3c�9������AGԃ�E�NJp���y��k����q %��vG�D'����"�y��ꟴ��� [��q~,v��Ӌ䭅�+��F��'>��_(Q�,����OyC���H([]�'6ѐg�����uǍ�a�z��r��h�������0�Y4��3 �����)��bSX�*��p9l ~&ꟐFl���6Ӿ���}PE���wꘝ�e����
ٮ.4u�8�N���d
t�^c6B�z�O�O���tKF�D�Z�q�՗����1-^��'���*�h�]D^4��γ Z�_�(�����xSs�'������H�ƧQ�^�أ�n���Fgc}�Sɢ�t��6�@�ƣ�y���Je���+N�<�k� (��o�l�[�"��F�ں��J#Y�:�ÊI������W؏0��U��oB����y���%��ML���%B��H=c����$8c*�R�����<�^�u�W�i�qK���ׂu��=a��}��F�f�����M�n"s6��ON?��Q,�G|���z��W��5Ś� ?��	��?���^=Ժ��F���(f��0�xTM���^�ת:�]RGơiC�[��ed@�����w��׾٠�|���,~NX{;��K<>��q	�=���/�+���F
q*s��~��snц��toS�٘]�_�1�q�qt=F��<����:[#l7�G���\���ʼ�'�;�����]B��f/�_.�9){?���m�q���>�B}��w�: �~�v��Ib�?#j�F��B�lͺ�Fקx���Kx��c6X՗V���J�5�H��UQ����v`S���;�*��e����CM���W���j	r��g< �|��v��\m��:$�;�a��>� Rο�⊑����-���/D ���Cq0��3R��K��B;(�ۑ}�jH4��TF����Y�0��$�b�Y�K՜�Z�V1,Þ�OD�*�}����F$n��dO��y?f0QԎ�A(K�qp�UA3��^JK���OK ?$�Ϥ������b��:h�7��/y���e��
0��o�[�r�L�C/�s�ф;��*��~K׷�I����QWH��R�!3�KT�L�uF���^�G4q/3K��G�Pe���g�4��J �"�-Y�<[<����B�ޥ7��lc臧?�JcU?�&Jw��g��̀®�8lóB���G��ʚe*���ng�9���h#<��S��2��@�Ś�����L+��:���̴W&�A���e�����\]U�}k��#:\������-o��)A���@\�ұs�ɲn��6����E��0�	2ve�����V5�D�TFՄ�Uݛ����AMڴ��.�^�x�q�.	��Ի�W����^3Yr�*W�L�R|�\����fjw�^�/����e|�V�r7hcܳ�jr��yg��|J����z�T`Kr�n@�>�$M�n��YJ��K�~c�Uk�e�rIh�:�����q>E�yg�(��y���L��$��*����X�nE!��o?���m����v�����M�岡R���C��7�Qw�����pH�"���s�v�Ѭ�R׵q�,?��6�X���9��	׻hI<�O�+��=�#�ġ��U�dE��AA;BXlxV65EB    fa00    2750i6,�
�U w��("`�<��Q�A@l��}3��I��鸳x?�힔8㟱,:�:�5����8Ɣ_�e}��N
�����	ev[}â�����=����r�-B��y�8��P�K��;�
�O���\��5���iıʷؙl��)[��Q������jϐ=�D�;О1�v�D�b�ķ34�]�8/��,�K�����;��׆�1o��P}P�S�Ƥ�^K�}�A�,F�&�l/��py�i��d�^ܓ1��Qoh��Ȩ�@���[&Lxy��Ec}��&�?���*p�5���-��"]�T��5P�b�g��3;Y��P� \�	��9ޏq������@�� �6�q@\���9r .��#؅�_汊nK0��k� W�}޺4�'�r@��@�
�;P׭{lu��A����A���q��q�Y��:�������D.�s�9zT��n뢊�������ڼ&t���̓5%�V�_A��a���uh#no��ԭZp�0��]�i���C�p/R�6_��!�F�ե.�����D#ۨI/��;��td�4�����g���S��\�ou\�������H4�.95����O%�l�P�+7A�gH,��E��aYJ���F���&���2��Oy��_��ܰ��*	+�h!�Fn�=����"��������O}��Ӣ��]8��"����]��2a�U5-c=�D�[c��q�K�w���������8���u�b*�^�ޙ���
b'jIYC�j�}}'N&��T�P�R���̜�W��wo�qD�)��`�z;Sf�<\u�`gz��$b���U�{Ĩw��}��X:	�~{������n������T)���5�>5��r\/&�?0�,I��/a������XC�炙K�;V�?�����Z��f�i�'����/�?u�ī ��d*�j�'3\�݀��0�+��~� ���
���`���tOM��
�\��-�V���@�i&ؤ�U5��g��Hy�u� mjyNz
U�`�\����<�Q����k76H�����x�	5��?�%}P�Ea�oE�r{�ز��ڈ��%��3�`�c��Mx�\!$��_Y G_{� �����R��ǖ�)uQ�x汪�V`y��d�#���`��g��]�D�|σ��/̘�����n�[�e��b��r���ȟ�֥� �VtF<j�JH�Xӛ�;d��<h�#Ӊ��{� �V8|�(��Fj\X��%��'�i�P���PV5�!xi��Q�p��D8bM�a����֑�:��E�͛ 1��Ƥ|�#�'��
_.�QE�#��e����j��?{ʮ|��g�p�e��&�BKu�,-�2�W��5߬�t67����	�[z���k>[���փ�OK��[���&�])h�=+����5>*/
�~��h�%y>��`�̛���)�o=������88�x��+Yrc�:�#v+^D1�����pF�^��<j��՘8O���S����.�ԯ6%w���|M�a��D�C�"]�������=�5�j���H�
i�8�h�����j@�������o�}�"<��t������)��
�T-ƌ��1�G7�|Ř�4{��D��T�w$}{���7��D��Ez���U�4h�����.	=���@P�U��ɓ%2�õ��Ƹ�@�+���q`
�#l����� ��M�B���N�!rN��=v�fNH:ѥf�����Q����F��)�\3J\-�T��V���EF��$����5Γ�	l�2�ؒ<q�p���Ì7��|N&at���2�~��,Woݼfi�j��kC���Yg�w�k��| 3]��Dn�B�Y��t�X*��R@H��Z�Ԃw=���h�������,s/�ΆH]�~ocY���d��E�X�6�JS+���ʈ�{�K'}��Ԑ�f��GiwB��V5	^�%&�-��ˠ�j���&*�C�Q0krơ`)?�@ 	�'��pu�Mՠ�˅&D������-��f t{j�D=RT��&����B�+a(\hfru���Ɛ��@i��hn3I5!:B����"M[�r)��\Uvq���Qh3FD�цO��N��L5���\�x�R� �����!�R.�� q�ĳ~����
2�|������U�3I��k�d����c�͂��F.z����#�ER1�(l�A���W�r�{�TE��{�V�VS!�X����� �wl#��#x���m���F^��N�fƸ('��ܹO?$>3���T�Mh�9���V^+w��NUL�%9�(�}�t�ѣf%���* hk2<���w� �N�� ��1E��h�A	�#�ԩo8�P�����.�/N]a)㛯@��N:���RY^�8=��m+��qZ>|��L��r�`9�k��� Vq����b��.�n��NXr�V�6(k�vi.�C%	��{e ����`4��7�cI��?�I)�5T�q���!����2����j��[�t�դ��h��5����:_��kQ�T�sji��-L~]c��K}��o>���7��v���8&�M��������F��Nhw@��h`Z�i243Ӄdd�r]��Cz�ݿ�{a�d��uJ4K8� 3��[��MaKV�q��0�^H��oRgng)p�LБ� ��Fg�b�����i$�RjzQx=h��ۇ]�����IRn)��.�#DoM��ka�[�;��O�4�	��������Tyv�ޡ��e�a����vzS�ϋA%�lhAl��cX�e������#5�5�.�2Ym�aP��U`uu��VKza�s� ��|���E�|V!p���J�E����?���hӕl@Ŏ�z�YDǅ�(���s��dM��Os��lV����u0�R���*2�{DC�؉f�B� /$���,�x��u�s(��D�U�Rf��  ���o���� �Y��^�����cG-.SG��]јon�Xy���Z)鼘P����	�~��񒳣-�z�kK��£Z�B2.�-3BO���m�ߘ��� � ��heXO��y��v��%�$ȸ`�,�����d	~<ܨ?�@	��zk~נ��:�Ԋ==���,�dF�|jE�J�|Dξ��g	wqʐx�<��g�՜r��>��ϝ�?��i!ڀ������)_������l@�$���A���a�_�(��F�d���T9��9�_�_��_Pj��}z�pU�8`��h֜v3!Td�oL߮�-��P��`0I~k\�2'S���DVn���jr���Pc�&(��1�\�	X���i�t��5<�GM�{�RD���;Q,[�i�k���cQ R;z*a����r=�Ͷo��^����Z��'�|r��5�ja�ƫ�<���L�h���u0��,�~�i�?����pz��?#�R���(��ZÈ���}_��]�X�V�.�#m�}*A^�)�j!�4��8V��N%����T�_[�>z�
/�T�iy�|y�6��\��ñ>7M�]������|�@�̩�c��KB:0s|RpWn��������B�'��$K댗le��Rbt�`��1wY�ds�uuny�$�l>�d�u����mgm�������2Q򪧳F�`9�:>)G�,�dCx�1���O�	Bm# �.�4u�v�x��x�@ � ���i[��J^�q��cqC.�H�JMg}mx)��䎶2G��$�Ꮂr]c�g7"�Ц���q�f�� Ŭ1[�3��X+�D�䢪��y_bx�~�&.HL�b��>^��f�!+<�9���	f��'øF�kƨ#����}��F���3�q#�<�+�ař�6��\:�*�&���`�9��T_�?YL_T5��w���x�w��x$���I�j�"�b2�7�r��U>F��N4����ۨOz	y)���߅/OxW�#���$����a�>����"�͉g[*���ӝ�<���N
S�ϵT9�;������;?��.W9�]%���I���R ���m>�����:��3n������VVZ*�vI����v*U�]g�q�
r���>�4(�	���s�>�Cg1]`*cklR�;�J�;s���|~�;� �Vzp��5��TXz��O�"FO]�YY�"qf��V�XCL�r��4�qSu��o���r����
Q�v��]�`(�����'�!.rFp�bwC���Y �E�ϭ�ъ_����B��ұ�\�9���:���:��b�Բ���&��8���-/TVԈ �W`��`�m�g��[��sۭ�ْ��!�T�&�S���!�v��{���[��j����{���eSÿ��D���ϭ\\+��bx�}�R�Q_E�Ղ��B��d2Vuk[@a�4��L�y2:e��Q�(�x`8!
��D�T ��E�f��Ϝ=��C�A2��8�ܑ����������m����l�+��`�	���k��X������si]ЉGYB@���"��8��>������~��u�Rb��Y�,t��F1b�P�֒�h��#�{���e.����^�RX5~
Y�-9�~M�
~�K��?K� P[Dy�bo��5�dR��{�^���pVeUӽ����Ė���X���	�f{�D�ƀl+�9����=��G�K<�$��~���D�̒�ܩׯxi�N��ł��rè�(���b�Ża����+!�v�3yf#�#�_oݚ6;
�z5"5���Fڤ�^�`^�f��6��7�=����ISN�mV���3�Ċ����亹w5�xoH�R�Q⑵c��eCƆ�d�
>�zf��A#l�d��DujQq�s�~�>�X����ʜpq�Z�/)��^�F�ԃQ�4����,'�]�{tk�/b/[��9.qf�#Kru^��5NĦ��FI���ݠ�;�)��+�F����!MS�skE�����R���lܶ��T�'{�5��:J��'�wR&A!�s[�����"�7�M����+j��,�MF�qzP� ���1�(��Nc��hE;�����р���Ipkdr�D��ok�8���Jwm�j�d2D�u��9�/���&����Kצ��p��~��@�*��n���7��;�|������%5�s�|��9W��Mҕ�]e۲XqX,i�3r5��3�o���%+:9�ӷ%y��c *��M�\��1�r(~���	j�L��a/�M�T��{(�˙E��G?�o���y�b���~��\7y�03���9h`�ɸ�X}i"_��%�[��ۂi?��o_z�)����.)��m���9&X҄}��'�HNbU�컖Q�n�N��Ġ݆�`*#��QP�c��rG�E��w�.�\=�U�w�W!Р�^ ?�v�|Y�ֻ�_��Ezb~���m������4ȷ)� 3�A�z����kjN֘^�Ц�y�e/��!�?,���Ia3�����l�A�~����͉�'�S/�JF���m��c���k̰^0��⑍)#��BG.:���%��a�hg�]���Q%f���������d��en
��/�s���b�m�x�ә�F��/�(W�p���_Xb��-��*�̚�y� �׿{v��<�O�Y������7���VPw:�3Ꚓj�-���E�D:�Ť�t~}t6��s����2�G�O��l�[ԃ�K��1N!��5�i�}�k��K�>�j��XՕ���/���e���no�fֶ<Ցw[_D
_T� ~*R�#+��X���MBv�x"?~ʐn ��g�_�����6��z,e eA�mst0/������AT/鬼!�.�t��V�l?�/�4��!td��ѦS�V�T1���OLo���W���~�|�i�d��Cp��Y�œ� �qvDJ�c���h�A�����-�ӱw5^�R�:�bt��4������o��/�=�jy��y��C���4C��̦T(;���ڄCe�;��Z��ndw������Jx�X/�{bhS��[g�b;��幻1D�W@oށӈ���!`ua�yz���~�t޻�*}��S���e ��� �����aK����u��ǅb���͠����b�0�i�F��0%}���h�?UQh�Fg�������Sq/�Q,�\v2S�iM��-z��ӳ��<���Q�he~%��d�d���.Ar�@����B����QQ��n����,Jw��B
�%Z4�/�2O�r(s�A�>���]42Z.$A�G]����3ْu��N�a�D�'�F�H9*F$}_R���=���1�A�coX�����8i���~*�p�����_�F�E/�#x�l����\��	�c�� �����-��a#���#K
��(A�ڱ�|�bG�m�����|��=f�If�2������YOh���~
�Ew�UW����q/u���ȍ�|
+%�� \9�����Kϭ|�aA�f�O�G�=ȕF疖&0x1��Ы��W���1��H9��:����+�[�{�[i��h�xr���ݨ���s�Ҕ�Ե'�X萣+��U�3��j�!K�{E�t��Ԏ���4^=�fA�ǰ\^�1�l�O�X���fx��PSg��C^��5U��WxcY�v��٨��ܐ�)J��I��E%S._Vt�	Fy��`��'U""6�^3~]	�����:�CQ�h�oz�����ִ��+}k�5?��Z`99ț��Vh���G*>7`*ʷG@J ����R��U��?��zn>a\� ����pn���]]�:;�H��(WS�� ^w(��L���cT�w��{:�cÄ��Z1�2*<��|��R�C^��f\?�3��b0�N̩-�en�	S�����-��12Be�"��V p��C����ǫ��#���e� ( ���KD�"�M�TƏ%�-�n�K�lA��.��X+�z-���CE�$�RM�����%�����?����,��;��'��U�^�6�h�դza)��'p~"q=!E��D�K�G����)s��k� ��?�c>�B9���,a��/�L�'��؜f�{2Sx2几7��4s`���G��P6@��>�$��ǎY-r�z�*��e+ȔH ~��P�b;�n�<��n�-���U�0�!���gU7�4�>�"�P�!����K����e�mq���Y�L	腷�ۼ��:���wn��U����F��q
!�u�5L#�����)N�tv ��N���):+6�c���2n!�ROHUW��~~�20-��s�]�+ΨrF��{~�v�~��=-�^��	�&���O��s�ц�?0�:�/���P'H���,{tx�S�z������W��ӊŽ�l�.o>L�����q���4��a�Ґi�w�d�
�@�@	�@�R�3����ɪ	�:n�q!P�d�0�vթ~`���k��h�����퐹h̏�5�U����\���(���P���fl62��@A����d�IуO����fX���6"���:>&UH�P�
�q�h{�;O��ߜ��xjŗRإ�������x�{&�d��^��Zb������d�Nֳ��̮��b���P�e�{!�����2_;C2ˈZЃ����V�i�=��$���l��w��ǡ�)��2[���(z�z�z�]�LkQ�Tr��*�4V�Mg�D�^pu[��`�{���I�*��1��m�5˶�K�L	 ���ƾ�Be�-Y���iJ�ާ�XV�h]�e9׏~v\}�u�淒V�=�P�⁦�y��3ec�qv��1,C�Rth�(�(�Kdy�h|�BK�Q�Bd���x�=�5U��=Q�>�=X����������%M:F?K�0�w'3�/_�W �����훠��q������z>03|��CJ�\��e�n)�r˲��J�ozD���d��9s�����U4a.���VN��x�Dq�	k.�u�'��ww���Tmn!%*�<��=e��V��y%���aSx��P���6Ҵ����o�^r��NZe�Gw�����NqN#����u��L��S*\"7���@L �뤉ݘ�A�p�o�?�,�]�3��C>*���T�Z�@w�A�6|�zs�@b<2�<�/h;�-91s��j�Sp�`s���������ד �|QHM�=CΝD�{�A�j����2���إX���u�U �v� ��Y@�E����dN_�`ט����6d�}�6=	e����%�8��f6 ������O~y���*�~?�Hr�\Q.`�N��B��$/Jq���t������ח��g4��><b����6�$\�ogÃ��}�`�������)��A�wW�X�=�����1��Ւi�t�lg½���%Mq�~;�C�tl�q}O�I�#p*�e~� �"6
X�'�mr�q���nY�����/�߱@R|������{B�Wz��+@�=��A� n��ʹG*�o�������7��	<p]�S��ۃ�fY�?>s�z��~^�|��:K'�#����J�9N< �~� k4[ �6*Hٙ�N��eo��>���@%UwPe�� ��ZP�=�I�x���W�`q4�u�b��Lz���N���f�N��h��g�nt�N*q� �{R[�?v���J�߻QF��[��F+�>ZJZ�%��]��s �
U��#��K�����_�#a�f�L�f=���{�BX��Py�u1ϠY����e������R�a�p��aׄ�R�;^��
�+tM]�`�U�!���?����`�g���6Z&G�ү3n��^�5Xj�����/Ӫ��~ގ+���^ePza"��ۺ��������C�8��
�]ҒÜ<[�ח���J3%�P-c�(�Ҥ{M�2���Ӎ���E����]_��}3�r��'z�\w�\H��R̒CIg�� �|�D��@3�_w��w�r�k1X����缪�O�/�Æc|M�.6��k#wE�+"�;T�n��b���;�0�}����Bc���7�h��ܵ��G� �'\5'��g���ꦏmQ��S|�qw�|�~���US��Sf�|��_{&2�K<�*4k�hŮ��oW���/���ɼKw䒢'AE�*��3� ������G����Ts�\���ҔO4��Ǎ�v_i$=͛m�V|D]z��(��u�}�`���?�>F��4cB�R`g�3%8.22yEh�� VAom��o�zTW��Bd�"QƽλG���!;��-�s�w��1�L�=x�0:���ul칎B��� L|�< ����^* ������zVt�W笕�̽�?x�M�9��I�܉N}���èB��z�<1a�yk�+�'�HH��z���cr��$��q8k��&Ǖ8F��6�`��T�N,p��6�B��rm��G�_��3H>F���%�n+��ڦF1����ܚ��;�>�y.gN�T'����-�4	>���k9=:�r�H��H����h��Uz�w-as�o<��)
��`�D#ΰǶ�͛�AkmUt��f#���~�`*�A�wh�<\�*?f�7!"F���X��Ǒ��k�#$ׇYpF�n�ٲ����L��\����G�2^z_S%rfeJB�� �-r|ԗ-4f3 ��Ů�C�|�D�_ѯ������i�M3���Ak	E��^�����|Wc�����l���R{$-�}�U%@���{������U�k���ƣuu��֪�/�z�W�6�tz-d�K���ô�>���Wd�H"�#�p[t����q㖊����D������T�6WWO	h$��{�z�o�6(v��2�M-e��2�I��3�<Q�v�cp6MB�"Ȼ�𴵍�&,>�2�l�q��>�"mJ��VP�Z�o�.��[�
�����v�v�l�(k���s$���u��V}��\Ϩ?S
.z�fµ�/��Zl�(���y��=-N�l�~��3�O��~�	�T~�K�"3dcn��G0�;��#8I�C������$b	=��tm m��:sXlxV65EB     2e4     150��3���؂�����|H?�������v��eI��5�b�	K]��l�T�>�'=n-�IN}�g�����V;�$>��dR��0	m�Sq�C`3n��q1�By�T������P�[x�Qi�0���X~�?-��5X�F����ǉ(������MoD���O�����.ȴ ���}�k�H|R��FtM4��'NT�R��U�N@A+O_T�SB��+y��&Ĉ�	�{���#�$u�_eK͖�st�0���l6�E�h�\2���N�}��KJ���V�����%]�A�(��گB5O��L\�j�ߑ7Jl�	��������r��\�Y�+�
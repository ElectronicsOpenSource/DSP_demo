XlxV65EB    325a     d50��M��"z]�t*���Ȃ��n��i<N��I}2��-�A_�?��LKy�$j,�>-���*�uQ�[u�d�[��R�<e�m��B�t{���>߅�l�l/n+��2���h#R �m� ?��C���)E�o���[�؛Ҟ�T���i@l~�8�b/����N�C��j$5؟�Ys�5�~4� ����T�b^��Z~L��AS�%˼Z��.G����s3����˫f��s>7�؋�+�&2ϸ����V}}����s�t���#��zֽ5���2��V�=����}�V�#�����ҝy�S����HO��2F���vo{
��B2�N�AH1�|fX���sL���d |�H��,6�;z	c	��Z��0���g`��7��Ċ���=��,��M�����I2�Gע5 KMq�����+�2O�����\��$W��ͱn9��Jp��P%�M��^`�C�	Sö�t�i��Y���ӁdL��Y	?���C��{�U�z�q�F�p�E���D[����L�����`b�\�F [ò¢"�6���E��	]z,Noxܷ0t� �U��֎��g��#��w��1h�2K�^n�ZO5%��%�v#d-}[�>��&`T�Q��.���̅W� Ӆ��S�T�0���;��k���+�ax-w��P{84��k�.+�x�
rλ���U9�魴�;_5�pI꩸�ڡƃ��ۙk���3`t�0ڸ&!W�Ԣ�����[�q���zb1�~>�WY|3�z��ڟ�N�9#���fx�jk>7�M�|m��l�		���O��z4a��q���t��s{�2^�%N�K���r�v�L�Y��Q&o�"L�� %����9A�M���V���N ����2��]�����84Fphh���	ݾ���N��8�S���0�������&a��7M(lѧ��w���j%���ĄYO�cXbr�7B����G�fE=��"����hV���%ڒ`��k��9A�o,bs�Pa^�z�.'�as�?}[�A	�D���]�Er.g@�݆O�4u~wytܣ�����:�<	����ܮ	����d�#>st�;���a����]�gJp�VXL��'o�m�Q̹R�E�R����
Si��v�:yی��ʮ�WF���("c5�~;�"@�<�0e�A�B��M�_{*�S<����(u�A�	8����/i}��W:��٭�㧊�\i��*�o��0[)H?K���;v�lW�֦��h����h�7K��.kܭΖ7}\8N�H�'ʶ�[�\�i��O���I�Pwgɦ8�Xϥ'}�A��r���Bɴ�#�{��%�O�vX8��
����z�M8`��+J���]>�AzkcQ���i�7n���1#�%����>�<�T�@���c+Փ�7�l Lͻ�=a<�4)���@@iE��2���{>������H������>���H�c,���Z��qc��|%~�Xx^ �.G[��g�4Mp0h\�1Ɂ�&�����8��`�S�d�\Ypp����&�:%f����k��{��b�3B�������W�z�#���Կ|f��� ���;�'8�,.��^�9���_����Q�ܲ
���ИTt*`ox�FtU�!�V�_��q���N���k���|G��ժ�,����>Sp��>M1���0��6�'q¿���h#ґ�S�ɋ#���*�[_�)X�p.��ns�}�>x5���]�/3�T��e���H�c[ʑ�2fhg?0Zb;p���eA�d/�2��t�4B�z	��m`Ӑ�ri�}�o:ia����ik��)�������Hʁ�Ñ����b���'D�a+Cߢ0���&�ظ'���*Zp�y��řh-��y���.�˻r+�7S�E���(�Cg{�Ĵ]��<\�9&��~ őF��:�OKΩ�;=SŰ��>�wb����K`�L��kݾ�.0��Fx�C�3�1mB�HBi��|�"��m�6��F�r+�dW�|?;��͊Z���8�#jK�gO�S�"o�`l�0�C��QS��t��=��W���,��I�vOb�e�:fܡQ�p's!!��O�0��ȱ�cQ�6b�%J#�*�ͪ)Z+�`��Xx����5������ɛ�92�4��O3�}�A�ԣ,Ң	>����B��V3�΅s�޻gc5d����q�Y��T[�y7��#]�Ys��C]�.�cv��o��i�~�ƴCnlI��]w����d�Q���b$��+� �R�p$��o�" l0N�2�$�2�v�N{�O�想�������15|����i�ε0�YU�)�g>3y<[N{�a�@,1b@�5�Z�}hr$�)�?��I�}��g0� q���Z7>f���Mkl|苰W=���VUjC�;؂u#���sX�5~9��>�ER�[��&�Ō�	�����6��1�٨�� [�����N
����#{I��7����g
RZ)�vn�v+�Ʌ ��x�<n����5���;P�z��7�̌8���º5��#|����xg���HMF	y�S$���2��Z�W5���KKa�'��\f�&��P�������x"�*�b�����XYw��t]�6�/�6'����p�����J�E���6xT��Ͷ��F9(����8�����O�$�&
ߊ�*���#��%��U�?�c �.��T&��$s."y6����z�\�>E�돭�.<q�KS�	�5EX���:�~�$ᮛ��\����`\�C��n�x�c����Y���!��3�Zk+�]��>���1��K��kZ�͘�, ��ԷE���f��!7����_����2M��_�Ņ����.W��+-؅��2	l@����ȡ����DS)�Ы��4B,�qv���m��ҫ^8��X���`\`_�◥S655���h����֙(�@��\7o�Ss��g�$�dƚ_G^9EjЊ�T��7����E��02}���Y8Al*�q���������<�A��@ 2u�S�C�kϥog4�r�=Q���^'$��g=�4���r_K��{�!3
n����vVJ��2E
��>,�j�Q��ѷ2��~>��yߡl	��tit�V�hǂχP���Z X��� 7�莘��� �1@*c�~EX��N[��[W�}h�HP�}��7����4��U'�3�Zw< ����+�qm��s��}LY�3���Ye���#C�1r)�$��L��
�%=qC2��`+G^�u{�aw!@ܸ[+�0��R�;��o�eXd9��[կs��b�*�l��KlI�;ꬭ�.��Pe���%�~g�j��>\�sr�O'�$.?�L M��uIS
XlxV65EB    198d     830���}�W�4I,'���h��<���vg�E"q��`,�8�PƹX�nNqo�	�v�.ԝ��5I��px�-ʀ@u�+�����3�Z�g� Y߻��\�����ֲ���1�@�վ��(� �p�cV�(�$�=����t�zl� �,�Pp��F:M�S�����_xkb|�t��)Є8��6H
�LW�Nt�Z��W,;��s0�q���\׫dD�MGT�Ҿf���MF��\��Kf�)�Bv�T
�F:�#)���,�CR9����dT"��p}lLދ0Z�ܲ���8�/�� $2~Vb��u�0��r�����@J�a����cB%>��L�p���	��[/���J6f�I�!3e�
X����GT�,�3ӊZ�����q��+_�l�D�S�����'T����s.���g�n	b1�M�N���I��b���W_㍯sӻ���ŏ�A>�yF�$��I�c�
�̸��9(�� �.��d*ϔ���n�LK~�|{�Z�=��p^�[:d4�[�<y'����Nꃚ7��Mb��f�1�Cd���d�.Hd7@ր��+��yIf�F�6Ȧzw��TF�6�%��F��[��ׁT�^5�WX�����w�bk|�!��C~Q� �k�R�5�|�u&��	>��u�pO�=M�`im�M�%
R��y5���|��z���w ���S9ˑϫJw�Uڛ�ֳ�`�B���vw��~����T�+��=�r[ڵ�?X/*!]��2a��,U*����E�@�6H0���j��JH�>�h�l���G�{si�U^}X����ʃS�F͡�Q.���F8��V����E9S?���X�R�)@�-@ߤ�����k�����[kx�q4Fo�������@&�U�����H��d�$��_!�K*1�k��U��Γԯ_��OF�Zׂ��C8�j4*!7�w���ݮf����>��~e�!� ��]�#�wTel�k�vF�i�[-@Bd�����;7A5B��@����{�/�8��{��GG˛:?.N�4�M/s��iڙ43"ZŠ�1���XU��fC����t\t��ݡw��d�(�W��;2�i�W)���c }L}���b�rId#5`�����o�*�@3h3�����ڈGO�}�"�d#�=ҸԴ˩>�L[�a�OκQ7ԓ6��0�� ��|�n��~�DY�q� ������6��u��圗�_R�7�U���!j�l�!��C��,I��kn�(�*��[��C�܋��˛�����t�󛎆�� �������w�s�#��*oqSs� �S�4}����(G��d_U ל���v���נ�Og���ɻ�x)��״�|;�j�E�j�L36��G�e������~Oh!4hS�]FlkC�P����r>��Czx�˛[����^��禷d�^T�c���X#�H1��/G��?M��r}̘}�BN��'�V"M�.�	Ϛ�����r�k��$�p�w�붔�įM�7N�:���(��P�O<��K>o�9�Һ�2<�h�#���𢡊��X2�ɂ7� 2L�˹���U%�Gw@c�����/6{�eI$��g�*�@j����Q�&�e��vS|�HX�����n�԰ٷ)Y�䞀?@5ε��$�5�$��vc�N!8�T3ͽ��,L!�.cdR��J����	ȋ��DΩ��	�(?D��L���-����M�jS��IK�5ù�Q�a�iT��I���ܜ.�HLx �/׼A�(?^���D0jL^B�2���
{U���6���x]ɹ���'�6��_��)���P7�$���}�� ��W�R�k��a��ƺ�QH@{3_����GT�۞��3-���������w|�VH� ͫO(����2nY���f���g
���
�L�0�J�������LC˷�N����y;���\�k���ck�嗉~���e5��. �E��]�ͽ���_�U�_5�E��U�/Ԯ�	��Ό�~��9a7Z��{�z�g7o��$oh�\�p�!�Y�\�,�oS��:q�xtMY��-_|�i�|���E=QI�F��.�Mh-+���nFћwR.X�J��a|
XlxV65EB    fa00    2ee0���M?��0��xC��L=i��"��{H1o��� �#�xa���-	�F<�\0|�����ٌdBb9�#�A_~I��+�(VIC������^����%u<h�=���5�H��7y?�?@���
s9a����К�;�BbPэGsG�~��B���b��h���=uo�@�*���?��	C C�d#9�z�����x�	������-�iՊ����կ�M�U��VW9$<|$�V�̨fZ,M�i���k=�����k[ Տڲ�,��,�� U�F2�����En��Y�B\�]�&CR�H���HJ|�1�l	��;���+�s�cu/��?���х����5�r�ʎ���?2���+F�,̄����7���(�9����6ZV��<ۚ�+��z*kM��w�l,>R	iK����/۝�N�0h#9Y����kqY6 �z]���~ ���Ӯ$f�:y��D>�C��B�{C[�\+)F-cQ@�̧E�i�Q���y"�64V���حo����H��v$�$ �ح��P�3�f��N�Q�^s�A&d,6��Nf��UE��H>y��dq~{�0�q',�H���.�K�p(B��t�`	l��W��5�4�A��G���V��b�-�|��_��u��xf�,�A�CU�:#��-cԷ�O�f�Mjc}���\>��\��p�4�#Ui4o�Ŗ*��,xS��IU�w���>��w	7��)x��;�,D�F��'6Gگ�`o��=��
:� t�ztrF�q}"2Oً��]	*G��#ԫ���ƈn���%]^g�I�:"�Ș^����H�)���eSjE��B���YEAaەZ��=��{����U=.���1w�r�O�+�1=~�����OF��>y���U�����l_g��[���,��_P�÷�܈,���\*:%�ŉ�g�]9���d؅GWt���nE	������k�%�a%�$E�hL��Ì���Kcd?t��z.w�Ҳ�Q���Q�@"��F�h/�S�IXh�B�Z��;�v��X��@Y�ĘWO�pe�E�%��U5L�ZPz�wsN����^CK7��m�~����� ~��%}^Hi�
���zȽB��l��ؐV.�х��LУ�lA����+�פ���mS��(�����{�E)�8�a�-A��]S=	�ڝ�-䇧�>�b�զӏ���?�G��?����~�����J��ɯ!�#������& ���Ud_�= j�f��������#��US��ȁ�N��sc��駈�qm�XNi�8���X����+���r-0؛�wO��E��P�K�ۘPЋoϻd�bԝ㷶��{J�&!���B��p�_$_~Iκ9יG;=K��I ���l�.Z�9�s?���B���g�
���!c���{"�����_���[���,b���Q�I�;Z�^y;[���y�KC|s�d�V��%�ݎZmC�[Z�Е�C�0ǐ�_`�{3#�|0��I��6�P+"��WC\űc�&qդ�Y{�y��\9�7ꎾ"�!�)%7Ǡ�Z�A�LL.�l��Y��^�8Ș<�����TN&���䓶G��ᾣ)'SV��T�vG8{�!��r��W�Y�I�z9*�[
|ec\Q�I�"S��"�G����g+ޒ�;��;3��>�8ؠ�)]�[h��}k&IM	0�XZ��F�t3��to#
Y+M�+�P]ɷ��a�h<}d��/�
\���aG���R�>T�`:1�e�)Z3�X����K=.�l�<[g����:r�ꘑ���TɁ|�RS���*��r��|��3b1DR3C@I%�+D����Q�� �1i��˕6��`Ǭ�'�V���1'����,$���18 ��T*Jv9
=��zÕ֭<��'9~S%|+��^��U��(��"�_�1I��2	�"ԗ���A�G��>,��N/��<j������j@����M%Si~��+ l�u�I��<��\�)j��s���W��I�R�s�����5+��Y��d����}�����ࡇ��5q�ߗ�L)K����iw���]{���~k��P�
�����`� �UP	�m�3{)A�����Ǆ(���]�-������p�%3Y�%�J�p��'����F/5!0�A�b�Iכ�;�Po��6�K�_w?��?*�&�ye_��)=�-p���F�5���,�.�O�1�������=fd�[�x�!E��D�᲍`�>�j�֣T��:�<��2&�)��ۃY6�¢OP�z��7���eF�t�����K�v�.��l����Jb��S��ݾ\P��#�~�W�h�s��7}S} ���-Tx�A�C�'��}�����-C�����V���ז�#o��(��s��)*��jy/�\�-��' g��X�z���[I���9h��KFB�sb6裴1Ò�����
��舜��}���6����HX&t-'\]X����٣�}Cs4i��K®�Lr)=3�bD��ld!����O�H�yN6߾��[gK$�s�)���Y���:�:C���Yy(�(<��E��)�$PKmYhRTu���J�i��I�f"á��s�J��(�]��<�+t��f�
����ܵhyWH�RW���RK�y`�.�"�ܤW���K8���JF>xC!M��.f�������(W�_�<8}�fI���d�l����Q�C��{<�`Vi׈8j̻�X"gF������8�4�����s_������Wp
�m��
����n�G֡�p��a���� �9�&�4\���?�h�O�.	�'4��=���>)7ڐ|��'�����C�)��H�)>2���Z0�#H#!����-��/p/����E	O� T�R��0|�5l�Uty��3o܌����eL��.��ǰ����O��d����!����~������;��$،�z}�>��{Hc���Q|ooζ��]���U"�ڮ�����3/K� $N�~ޏ�=�+�XjW>p��>%�~�x�������O�HTH�I����[�����<v�wJ�j������}�3��Q����7��������� ����r=m�[D�`�O/�"��6�ƚ�`l	d��
�){$�T��iӇ[��&1W����9�fG�
f���Gų��Tǀ��p�0l>�%6f�˘l�!��"3����������i���+��&��4�+:q�xɄ��X�Rj,dB�^�4���]��q�(G��.O`�@'�167�n�]Q��O.��V:z�*���~��ћ��Ζ([tF���'��Aܮ�c�[w��+�������ǔ��|��K Հ�?�x�nFȳcV=�+CFva[8��L�b������N2�a*�c�SW�U�	�~�67��2�g�e���#�LF�:���"�j�� ?)��[�Vo%`xsQ;J~e��d��`W3^W)|����q&��T�<T��#���Z��ip<f��������kD���`���gi]�I_�6�ҐD�ʕ��'ě��[�u�\~5���� ����b��{����Dг��������o����>\�Ğ�������ǆ,J�P�g�q�f���$lb���g/��4���eS>��&X�T��t�tu��91xP��u]�v����'��vP�_~�X��LQ�1����K_˩����>}�vL-�mi��Io�σ��E.�qIT�1��^����dA�%R�v+{�S����ġ@��Ї+����g�W�>S�X$Ŏ���,Crzt}�:�A~�#Y	�`����#������~46�=�OH�Z6�ۿ�~��[W|�f�{���-�mŀH=76���y`B&�W�ͷ(��T����E�u:c�H���$ꁴ�cђ����*����;�s�w
���`���w�8Q�Վ�)�L$d>�@�����k������&��t��OxA��}�����������#���9  _�D=H��B&,(���teb�ŁJҁvp�&>2b+��<�^���dEj.�{
Md�K�7g���e�M�t�}�A>-8-a�Rs�Q
��ڼ�<h�2�A0�b�ب�V�5�]t����̃ҙ֖��ă�R��P���Z,�VT6�h�:�؝��`�(c�k�gQ!/�e�-cP{�ɞ�ΘD!h�CR!��c���M/�����L�+�lI�ݾ� @D3��>c�?�ٖa2�G�h0�]�u.�O���1h$"Z.G�����Zѣ-5)4���N������Hts��	�=�r��/��S|��j)�
<�`\l!�ξ����I��agX�U�g\�TP�㘃!�+5��}����#Sk��V����C�;o�3���)���5n ��e��2�&�~P�mx��3D�7�w7�����$���/�KOj�r�;ãF��m3o-K�)Xo��m��i��0�h�n�x}i p{�[w�]�T���CaV)�]�����К~@���l�'x�4m���v���&a�:����_uxEC�_��]���f'�`�-Zq��O5Ʌބ�[sF�c����)��?Boz��"�6`�k�A!ݛ�^���a?;-J��{�}�� ���('�
�ʱ�o��������	,����=JBlfM��5�r��ZW�Gt��%-D���R��Mߦl_i��v�3��� ���0Xۄ�;� <=��6���
�I�E2� 4dH�ʟ�4��"k�or7�<F��-�6"}0X_|B����M�ۨ�ѶWY���ѣ��TZ(8w��:��\���p>�; ���ʏ���[|т	� �#�Mc!����*@� �fU��;Z�(,��3��.�L	]�c�H�l,ү&_�ͦχ�(��yw�{�uq~�ۻ^�ۛ�;����c�����^�r���/&��1�{�GS�yi.qj�����o����|�4=9�8����,���AlУs*V������+���(�����~��-���yߦW%��E��)�j/���%�k�
?	-�(u�����,.ң����0���!�߳$\��$�#(z'��� :I]�^��jj̟c�w?�o�����?���*d�WE唿	=�鉸!9�����+
 *\B�JXk�o��Y;v|�2��q�{I���y	n^ں,C�m;U�f�G���}Q�v�|P�cua��SӋW���|>�q�q̙�L��-,7QW<ԭ�,
����Ic8�JԺ"º��=���H�L��<%+�W��Hp
��K�~��=�����i��Fy�^r^�\��<��o��~�7:ѫ��\Y���0�2A(�ei�v��C��Y���ƀFFe�n����k��ztt�&�Q��&�YU��;B�7�����ͻ)���Tg0�\��������ޕ�*05���Sf���M���� \�n�*B�0G�բ�_w`�ڥ���ƌ�i�ĞaȂXc-��N����_X�sh��%��o��bS�o����LUI6�k-~�l���v�I�͇v:R�r�*��2Wpuh\ jzRE�&}��~�U�13�\�#���oSK�+�5�	>��"L�bQųfa����Ͱ!=.���{SI@H��}{)�#�M5Ԡ�;m�R ��	�9�̭2����꩚+���3B�&���a.D�U�n�X��#-i�T��������y���{�mV��cO��[�k�o#�*!B��B�K�r]u0���e�'�	�̱�9�=�-��h"e܁q���P�a�`�]�I�vw\F��c�r�P�)�yC�V�WG��"���CU���:r.������_�Qti��!`@���f�g�v�p?U?s���jCg�J��E��l�w�OOM�:�,#�F+�g;�쵚�1�����}o��X�J���nj�:��N��K3C#�(&����2������ ����6rCx�Y���=�?���D!K5c���-e�^\���+P�䅴������rJ�_�bjڣ�O4t�W�g���/���J#�i�ּ�a�Og�a�����l2�2����B���~�"b�wX��?e�b�pt������z�گ�VDf;�8�Aw|�S���*8^��(��D[��va�R/��U%��&Fo�2S8��o7�#�|�@/�8�=�`�E�V�B2�����y|*���g�8��C��^��]�Q�Zx�U�7�4H��B��'5ɽ4����_N��,-�q!�55�Q��n����E���q�	:х�P�l�P�+���ώo\�.�YAáFc��^VP�Уm����8�3�x\��H���=c�Yz�������P0 ��<6��ێ��Ժ�BaX����<	o;����6�T�Z��ei6�u9�k�#�X��1}���ř�(�߹��%�#�f��N:���f@�l��So�Y<�z}`���!b�Q�`��MJ]-8L6f�\)��<�>(��'�l�]	��ub��T%^�,��_��xd93��;@7�]�Lj�,e���Vyd�@�D80�ԣ倿�2T�.�HW�;7�τ��X������nnkYƉ��r���/��D�(PK�,�r�[>:��q~DƠ��]U����8{K1��l�7���vYFVNh�;���9�������?��8�X)?�XT	����м����u��1EK���w�-�t�35�L�|�RJ�#?i�>�F���V��F��X�h�'6�L���Bt��%�������K�S�4,z�t����^�a�O��<���qtV���$�B���Uh~ѝI��vŰZA���X�_��@�`1t�Nmp7��oVd����X4ԓ*r�:镰	<C�a�����Dv�%~����d9bm������|� 3ϰV<�Ϩ#,�kzi�M�y��T�uJ�k��j@f���˯~M���󶽗�i�j�4�^|��]mP�u)iv[���Oi���1� ;�g�2�*�Aij��ƭ^�pv����W���N ;}Gg��w[�jj[Vۑ\�\ ��B�E�'���UʐH�^�%���m�i��{Aio��\�ߠ���%�.�f��7*��X���G>��.$�4�E�s!�f��u��x��;o:��si�Cz��˪�w��1�'	��9�"�n�k���ֈ^�*��S%8������vں鷽�>u Z�=��i�y�i��Q�^�'#O��U���*G܊�XY�ŗ�i����d�;/�6�f{��IhS2��.���/*9b�ۦM6[�����ͷ�؟a��[��9�m�,n�j�'��flkCj�v��o�� 3>�j>�b�-�5hQ�Ø+���U�r4�#���k�yf#���)��?T���� ��Jy����9�w�����=�4���~�`�]�5�Ӑ�=��_���z�N���]�y�/6��-��#��$�B
�t<엧�[yigx���<��+r"�NV�伭%�㑀���F����3����v����1��G�\���F�p���v�_ZD1�,�\٨t��w��M�1�U��5�(��J�'/;x.q��P�a����1}B�k����t>��	r�Ұ�t)���v����;Ȣ��s������>�ͭQ ܬ�W╜)�\,���T���u*jR���*���A猲<��I8�Il�B}?_Z�d��Nǝ]>���=�)�����t�2��{ͅ>q/u���.(=gGT������ͽIm#s���< ��˖&��ں�҅�{��B2U�w�����F��`J���j�����`� ��m,��D=���(��ş�|��<9��_{l��@�U��MC�k3W@��>�,?_7\&�Vv4�Z��#:-L%�|��i\a�(���T���Ϡu����1�q�@�K�Q�l�RE'����U�p����o.���^���]��R_.���'�.+�&� k�%+��/7�sN�u�
j�jb�k���
�>��onC<��o$4}~P�w}k�[�S�d`��v���`X_���y((�A;�Ǜ�!�|z �B�i�2��̦��:bM<L��&>MdE��^F���v��bޤښ��$T��WO�T��Tl|��w�����y���)�2�n�O畨j�3I��-*a�\j����H�O�M�j�����ge��hU��:�'���/D�pז��" g��pF�R��]�z�Y(�"E���u|V�B`����cƕjމЌ��^���@�����%q���}o����0�(�h^���H�����E�������lyd��:�K��Ч��WՃ�	gˡ�:�jw �Ws���K9���:�<K/?��R�)EE]�:��j*(��p�:�jU��ͮ�l�@�v�ӑ�R���~u��p���-��2���:�~��s�
��T�p�	���0��9���v: ��%I���,)�n���Vpcr�;w�c���8IJ����U��������T�o��&�H�����ϗF�3ν�gw�^��>��w ��R^�&)���t������mё=��&���8��1�+�&8S�Z�s�:�g�/�q���>��Y�1m�����`ne}jB#f{H<��H�T�ڭv���M\�{uL^yEg����K�e�O�zx�x��݉h�{,6��a!$2��=e���]-8�7�N{&n���\����D��Yi��\����%dS]���ȋ����7d���C�B�h����Yu�r!�ݠ;��O��Uq�\�ف�oZ��'&lM�3&���MG�#w5�|g/�0W>�q�G��PM��k��R�L����	�!EU�Z꨽��,����6�݈���MB~1s��<B� F�\��h��E�(Y�
�>y�y�	PZ,�D�f�DY�y�[{>���Y:�h��pB�«>�ǷQG@��q����Le�X����Z�� �o�Y^�����z�� ��Ӱ��-�
Wޟg� ��Ъ�?B��] �S�O�;տ
APf&��	�i+T� �����B3�,�\�b9��=�wS@?�~C*0�!�[�����A�ba��Ƭ�TQ�H�A%�RP<x4θ-����c]�!�o�!q	��*��^�~�F�l������n�<����]�#Kx��/�tZ� �[w�|�ύ��>@u��=l�.�(�����%�a�j��ʴ5�����Zu�ė�bY�����/�����o2B*.E"X�2x8@����,�U�l�C<07��E,��L�T{�r+Վ1a]�f�q) ̸fif�¿2Q|�3�T��4}���Y׏b;�xw ����,m[� �v\4,Bب��Ě�T%��kMY�8�;���;ZZ�Xܒm'��ǀ�6�-m���a0q�6R�_NP�w�&��
�^���~�%w,�aÚ{���/�e��U�9nY�9��Q�#��1C�GO����ً ?�/�u@��.�ɶUZ�_"n
zd VUv���CL��jZt�֊��oIZ�\�o��E`�r�Wo ��p�;�m/�4���"8ed���y� ���>��O�f<d���?�N�zPS�h �u�L���a^���4���������!�d�\A\KV�'�2�~ y��=�tr�2�yH�P@V\vFGƑ8�:�ӉkN"�d�\���B.Qv��ֱZ�c&����U|�?|i~¿����R3/�$ќ R5Y^3ͳ�Z����i����x�9y��g ��&�]�xx�p_L�=�����wf���o&!��X��	LI2
3�D��{����c�>��ەy���Գ�=]w��#����|Fh���!h�����j�N�Vp&Rj7(�A�adJp(5��6�����N�7�ٜX:u�~*fQf�;�ܱA�{�0�Jy_�zoZx�4-�諣	]m�\��Z��3OpA�%�»�f�O�>I��9�\'�A�5�ͫiN.vqO��!`�~�='�-�#�.��"�����p=a��2�q`P*�V�Ug�n���7������|8d�u��Ւݚ7?4�#�pK���#H�EC���)�"������@��v��y7�;^�BH��Ԓr�,�M��[��̓����.�R[�k��>���m�U|j����3c;F���pwfB����q������V���89�����xZ��G�K�'��ȅ�q�7�fq�_�~b׻ d��3��ѹ�L��Z\J�R�������t`)�8�h�j�8����o�C��#�x�s���r���$I]��T�l�����σ�7�Ɍ���V-�|;�u�RZ�\��8��@� aSCes0�/X�]�~���H��\r�������:��eSF�ؘF`�u�&�{0�m_�\n�05^��uB�rh$Yۑ >����hz}���0�4�5V��8����ƒ��ە"��#�8�����O�P7>%�Q�<���w�����̛b~A���gT��8�S�������KyC��7Fl�u�<�����mw�Ͱ�%�dEWR�\�X�D���T�4&	M���@2I�b�0��t��<��,���蚸	j�ڑV���/�w7BB2v�%�uB� �"#���O�A`���͋���� ��yO�(�D��r����`AU�̂�Nt�Ӏ����Vr���%�3�U�x�ĽѶ�� �4�o�c
�a9��s��X�#����.iyI��gT��k׭���"��E�|Ζp�X<Ey��u���~�ӟ~�="��g�E>K���~�[T ��}a�ֈ���B�l �q��g܀>[����=�;�O��QVNfKU/V��5C;�5VNvVT��_w��<_ڎQ���� ��h�Bs�4��,��f�Wr�݁���_}5�@4}ߖ&$�OeZ�1t������{$#/D�\�Ͷ��v������Zc��CRBJ������Գu����Ù��ٯ���,����dʃ:�7�R��y �I�����+(Lx���XN^�2T�r./L_=:��N�u��A�����D���j�|����J��w�\��uў��u��C��.k�s��n�����d�R��������:�Sz����Q����p���JtVW�ynnM��RC/�n��u\�$��d�W`���G��dG���;��Q��W7� ���Y�^�A�=%��8�K4 Q�E'G� �uO���j���J�,�4X�a�� ��J~Y���Rx���ְ�p���
����]p./��B�3�s��Z�9�ch�_�r��~��n�A��\�,�~�L�Ǳ��9��+��R��P�n��_T�Aؕ«�a^��`A�q�J�֭4&�3+��f��+��Э+ǘ�յO�~"w�{�H���15�qfԝXC��Xo���Ҏ'�����[23�r~d��������Q6S�W��(&������(����1�,�Ћ������9R�U/��g��4��;D��J���߶�p�6��j�(���U�z#�l兙�hk���*�d˷�@B\8ăe�Q��?�,��	n�bȄ�k�p1��;FQ�s��f�,�Q�f"j1/�I���1@^;�QXV�4�v��MoJ)\�Pⶾ��\��>]���^��j����L]��ҵ�5����~�GȢ��Q�2S�A�<�x�L�m��C�o3�Mk4A��x9��Z��`��������֬�y	��IZmld�p�p������-L�jG�f{�����z(Ç�:��A�* �p��B�v�'��o���AGD����ˣ�y*���'�壄�H[]TV��Q1�� e�2��A� ��|���Q��(fZ�����2�D�5��E������Jx�e~\Rz\�:;��(&���Bjs�'�j9S����G!��;{�rB�XlxV65EB    8d9e    1910-��;P[������xy��1z,;bdݝ�z&r�E?��*��(�E��/A׺�ҁԴ�ɯ��2�\(���7�ZI03��rÏ͹<���d�x:����Z5���>�kAћ������Js���O왎��bhfSr��f�����X�����D�"GW�*�ɑ�,����,C:��yK��v�`���Q<q&����\�����Nr��ÙK�#�+��)��Me�\L�c(ɺ]z�l��������UQ�ۗ1�Q{���5�=R�XB��ڤ�?�U�,ZU�28=П�uMs8y�� #ЙBu����3��b¿�g#�.��X
�!1T������)]S���_Q��z�}G,��q�����;5�wzf�!������tL)S��jT��:��#��~6Ȇ�����?���y���+�%�iV�;(,y� x(ϒ�O�z<�
�Ӑ�i�.�\�6S���(����q��jW랯$<�)���a9�|>?F�=����4P�J�d�ͲU��#I�Ȅ�v�
b�b�"/P.�JC�� &E�rET�i��^\,l�e�O?���|��l��܏Lm�"8��-�LF�3H*֣��#+Pk�����a�OrVD�\��+�H�ߌ���<G[�8���
M��6$(~���0��e�����>��h����hp��S���5_��q{����°��D�c�/v������uS�=�B�jy�Uok'r��$�=��P�1Q���Z���\�&J7pS�;'D!�"���#3�ĉ�B�4f�R���)J`�\�K�u~C�ah(��k��QE�`�CGW�F�͆I0g�S{;ޑ\�/����&������`����oՌ����6�2Zۘ�[���I�}��IY���F#Ɏ�> ���|z��X	�(^�����m�g�;�g�y]��ԌFeݒ�����n���`��Ӏi�Q����!��x�N��"�Y��{�퀍E���Cs�N��x T��L	́�F�Wj�rf���P�󋨖+V���g)�������6N���	���!��~���!RE�iO\�V�p˼U]f������a�:����=�������7�E#f:oɒWrw�ÚB�;.�^���s�#
C�`H�(o��~�z�� ���4u������W_2�����$(�F�O��}hf&[�s�*���dE���`�]HKs��Fl�����Vd댳�ɋ�{Z�[Q-7�VTb �Zƍ!��b��໹.��Z@�o�!F	��^�4֞ԋ{���l��4~�?�4l9��i`tY������1�#��x� �R��õ�c�1�q�F@���qnPM��ƿ�#�G��&IA(���;ظAsJ������L[�Ń	�\#��>(@4���~�+\�[	�%H �؍u��;�?f��e�薟c���)��:�k�s� \�C���	I;���Q"j��#-���F+�A`�X�PP�����]ގ��s ?��߫�I]�;,ۢ�|1ڋ�c�6������V�����%�?���!���+B�(Z k]�P��+e�
�b'D!m\0�Nfw?,`�5��I�;:���v ��Y��/17e��I���y@|Ѥ�	ݍX�[��x�f�Tx��j�"@�T���2ͬB������ֿK	�9�M:������ |?�:�k���_��ݞ���J�
����V̜��L��s*���:��/:)�f��
�Ay���Πʘ_�&=����������ߐ�{����ɲQ=��;�]������.>q?=� ⫵Mi���,���ӂ<�|~4�P�N{V��14�P'��d�;uZ�SS�Y�W�:�������Tk�uf.�P��]nBǂ��pc��F�eتZ��G�L�%?�OMm�8�#6	�$�?2B�ųH�m�qc<�A�5alpt$��k]c8<���vm|&c�V�R!�Y����g�l�/������E(���[�x�g�H2�i��^p�T-��kh.��
�-%�B����F k%n��Pґ��)�|�َ����zZ��M��_e:�a1�	�>�
)���Χ]`����K��Bউ�C���0�\�R�{?�o�8�ЗP�asTD���>�}�x2\���������K����C� ���J�v����$�r�$���/z� b6�jM�l�SR�ɺ���|�����#����8���n��	���^u�\B��3Rٖ{�7�<9a;Cy/,f�<�n4����� ������5���DL��3IQ�^M�̻������]�e>s�aPo)��q�aoj"٥}y-))c��;�,_�_��HX��@L�J����	T�H]QSՙ�ūR��C8a���ʪ���-�-�ޜaO!��|��'��p3a>�\6��t��e6�l*�Nzk����x
������"%u��u"�����A�u�`�xP'���\��@?(D��*7V�Gz�W�~��[�;gA�$���?�P�mB�<C�uɇ�q�*2�.���\x��!��1�.�Jk��ă��\�Og����$.OR3B�l��@;�F�o��������D�����9�a��s�_��s�>�7�KK���0�Ҋ��X �us�]�k��|+����/�TY���P�C�2���ȉԵb
�������O]nEJ�&g0g��H��n�I�@��z���.>R�,���8A��<�	�W0��쪣��{���K�؋]��s�y�kf @L6�P���3`B��X���uX��Q����~v,/3�K���z5	����1��F�q��S�,����?�<��P�hvkF2.$L8Ҽ�
�VF���I��/
M�ݳ��m��4�1߃�,�[dL6@oa�*�>�i�G��x��$�U�@�*^�e%^g�q��r_G�ͤ&M7�K�w��`�k�W��Gt��4�f��|o����#�Iv_��R��:�Fӄ���m*�zh��ۏ?d7W(N�d������8 e�A�ӷZ�C�gڻ~4��8�#��
�=�_�5��Q|�A7�ܦ#������识����U�Vf��w��.�.��x��G�/u�{Y�a��`�fx}_���� w��~�D2��Y;��ςsy(MpK�0�X����lKi�B�#�z^����Q���	]1�����TW�e�%{���/�V�4\�CIT3v=:\�\�I�9H��=x}�ތ�'��+��W�1XHH_ݗ�ڝ<��H��2�zɤ�@����`����R_��D�a��j7`�s=��~C	y� c�B}���5��#�������j�3G��lCK�$M�m�,�ظX�ϋ3�u����ǿخ��z�|���rB}s��l���}K��:��[����FP=;[j�[�:�ԧW����.s)��>�8ɸ�(뀊�`AN����O4Aj_�Y(�̲A#T�w.?ʖ�[�G�O�hw��)'��	�X-=�D��U�JcW�"Q_�X��(/�9z?���䟭r3nH�?Jۣ����|����+1�h�7{��k��ϮR���r�1�ݶ~��p i3P<�e�#L�&R$u�Io��4�*ی���m�+E!j=Jf��b�*����N�̲Wxc`��bڍ�rN���`�ƅ��x���,S�bRl�*ش	�|�e9.��e����n��pC�F�o�|��{���>�̯б8����b�[ ��ae.��#vפ��$�Y���*��'.�޿s�{�t��Xq�w5�d���*P>��&��U�c���x���N����H.M�<o�`�F�5�U�a���d����m=���0���V)�U�9�� ����RY��w7&w4����#��aj����r2��^LRXa��X�@��oQ��pP���Y���C
}D��g�d���}��>�����(ߡDX�>�Ͳ�>��B QK�VVs�7"U�nԼ�$�����>�x�0]�['��2 `����q�U��gh*6��5�.��6R�
�&���>�d�����W�%O~^tpI�U��0y�z=�E��(Mwr
��	�F�.��W��[���)ɠ��+=ECfl4�>
uْ"K�ɤ��R|�Xk5�N�?�ـ\��*Gv��L�yIE�756s���:v�Z8V��p\iW�#���O�J ���(���PԐ�]����p���ũL(�gI=����D�K��~h:o�{���clPY�-�L+�9�WV���(�a���t�b�Y_��܀�KOH�c��\�*��\�@S�1D�A0~�+� �Z�!&ۋ�:M�(H F7���&�Y_��B��lOAz�[�㧅Af�՞�u��J����E�_\G�}�߅y˰��[�j���`4��m�hm��t�2�9�@��E0ilg�ܴ��3���L�Kbb\����c���BN^��4!	l� ��U��lG�>���HR6�x�B������� z0��5):+7�/R�Tb��#����r~�eb�՗t�`��[Y#{y0���1[o�6���6H�8Ï���/3��?����c%��jKP����-�O�%�gg��.)���G�LavJ��h3".KՉ���ߧ��D4�n3��.�Q���� c<Z;�\M���nqjZ��	�/��W���8�wF�b�b:Y��/.N�"��yz!f4�����l�~�QV�����"��5ڢ�M~8uPwk?Sk�� ��"=@t@��oC ?�"�C!�̇�	��Kv����c5��h����s޽�-�����W�#���@�*j���l�N����'�����m*�Q�0�#)Y�r��,��G��)�%]��y7�������R�O�\_���>�v"@EQ.���EU�c�޼8TR�8A"�+�l��C>;�.���I���
�z�M�Ev`�3ԥ�/y��LJ{���O;?�L@�䁽ż��q�N9�X/u0q!���;'&J?� �ry-A�.O$[B!d�Ϟ.��y��_�|և����w�ѽ2J��,'��u"�gJ���)vD� ���D9I��e�s�GZ�L����a�k���"U���wi�^߿5*����a���~����l�`S�4����5t�>c�Km��ٲ:Av?��+ͺ����Ú�u��8ky��}($���Y2<��۸P�P��g�XH�^�%�-k��\���w���#(�s1��p+����i^IHWϾ�����W��^U��>� �f�}��\���ƾ��w�@¥��]���]�Mۭ���P�'&0����d��-�(�ɲ���+\v�O���W�7�Y* C�qml�c��da���ods����&G�J�̅��?!���*h	��]5S0e���M=�-3��V� �c�m�������%)��a	�A(���jY)_u�>�E�Sރ�|�YyL����Vk�i�Ţz �mJ��Q��k*��'2 _����_(*Es\�OY��=���^u��=������x���B���(�o!5m��,(��-l�PH	ƽ<��G��`^��J[WI���Ӛ;Sou[��]�?�Ϗ�H�P�U��P�܃���hu��P�OV,7��'�RDgg�Xt�I�b�c;b�@�89�$Z�	���2"%��a��-�z	!�W�пD�/l�oݙO�`{X#�qE�U_�ӂ�����h��ȭ�J���6�d�9X����3u�E�f.��a���|�D���$N�GWL�"��T6��:�t�]��??G�\pJS��PiΫ5��Y�F�`&Z�Ԋ49�1��z�(�`�妅i|���MMt�����ъ{�t-�ɛ�*dV׋6"�fˁ�n`�/��E����N���;:������~Է=P���3����P���x�-{H�2�i�i�t��2��3�kҟAā2��S�*wM�IZCZ��h������|��?�k%�M+C�E���M��C�:[���E�_xG������`���@j�.���\���UZ��5�}�pƔd�t���=1g��O����x�vc]N�a��_0����;�hWsҥ·�W�V��z�N�.�5 ��>*֛E��*�#,!�w���ķ��!����l��ߥ�6R�ss��
�L���� �q�Ό�2lv�W����9����Ok�H��~����A ���b�(_�-��Ϝ?˨ʒ_X�u������<��)�0���5�+��m溪^g,g.�-k����uz�M����r}���w���鲽�Ӹ��pwTu��+>8��Q ��TWW��ٶ2o��
XlxV65EB    fa00    2cd0���;v�dE`@+S)Y;�R�������+��d�4��\��8�,���y�u���
�N/_|c���[��XҖ�����	=Z�R�����,�ى�*��`"����g�F�6��N�[/�@$���I�+!���A R��DFf
�b�?����Sә*�T^e�Y��9�m��WgQ��g�-Ґ�I���������EA�-u�2bM@�*B�:�db�o�0�ɩʘ���4G����k�T��'�*�+հHΠ���י�!K��(���T�چ]�x��K{�).�ԭ�%q�2urzZ�I;�H~�Af)j��y��z�8�"'O�H+��JM&�A4qN�d�]���.�s=5�"%w��*�O��4��1��92��t^�(��я	6s������t�Ϡ��G��y��l�p�؆z�*r�+�B����ɵ|�"q�� 6�8=)�ݜ��)  ���{��{��`�j#8\Ħ|�xX>#x]a_��Ѷ��䅆�BI��£���yT�<��xo�7���:�m���Ex���4��@K�x	v$#O���DԆ�`�VP����]?�Y��U��d�8$	�H�+]ia�8�R��;%C��+�.i&�{���1�1�Қ	^���?����.��y�t�"n��ځ���|$�&N=�2;~
���]��Q�(EE/��n����z\�c�_k	_�S:,R�m�����C�_�Q~����X�hj��~�R�C5F�F����L�ޙʏ�@�z�Ty����3p��n.�n�kӖ���_��	�^[�0 %��4-�AT(�Lw��M0^G7u�m��T8���C�b�� �%��/>	����c�V9r��Ye@rɎ�`E\�8W�~�7�*��@���+��I�[�@������(�$ނ��p|� ��[���q���D��)�\�"<r یN�&�B�l�f�&�����I��D7�p.K�A�#�G� \�!v���hbFk�>G�:��H# �#��eI�� 6ө���?��=���߯˸���\3u{J(]�DO�Ƞ��:T�+�qid=�=%�o�u���Aŝ.�ơIE)*� j��X�6����xN��J;K5o���M(�V�Q�8��:�v)�⫝̸�M���"�������,�18�A�3�)ܡyĜX��������+�2
�����3�Dx�;NZ��=�+���v��x�B���?*
�ch�1nE"���	���vF�a\ �[��Ϫ�=����L�����򵔒?��eRQ�6`tj�|v?�enB��ҕ�8�]VdR @��'��>���w����+v�i����r�d2��3K��+r�E�7�X��݆���(X8��¬�A�����Շ]@�</�|`�#��$<9 H�z@
�Rf��8�,P'l�D�� ��W^���Π���:�Α�3<��NK�b��m�Kp5}�q	P�78�E�Odi���|���]��˗��򬈳��̦i���Y����Ғ���L홎��f(�� �cz:Y�F��pމ�n ��X�OH� 1�t���V�k�n�2m�CW��SL�N��c��M����BV��!'Q��G�sz3����EP��f��z*��e� ;'~6�'[��-�ι����tl^j�C�A���n^�k��MuO��_��yw�E�4?�,�]������e�w"~C�"mZ����$���~�]��X�raD�`��w;�{:�`���c���#���?�������K���2�:�II�s�B��4�����jX�p�IbP��Y ���/���B
"�n�a�0E/�y���s�%�b}��'�{��M�	"���Е��B�K�����b!���b:~z���T���P� " nL���2����V��19�^	2j��m��iu����+e7p��G�e��aZv\rQ���7�ڽ���ұ�P�aЭJ���������l��8�M��)%� ����<��0��e��5���h�A����q�Q��}��vē�o-+mG#�� �!��%<��G�nH=���Q�7��F`����^R�'ɗL��ܪ����w�tQ�-���mL��J8� z���K�?�ܬaN�IķPAr�<�2�t�}�s����J�B\C|�(F�����D���g'"Ǯ3M����5ؗ�)~�&r<xL"U�t�c
Frz�� O<Ӎ�s3$���-�w6�털�K<6�U)�<K'�s:4>�v30�֓�^�3**�����_�XJn`k�	���$�RC[�>�5�1���_���%��u�
:LX9�L)����e��"Ço�V��	P���������8b���*�Ժ��Y�j� ��G�ݣO��T��Pܭ�}~��֥4��D��^_9�*��aY~�Q",L���kLK���@;�l�a* ����e�u�O�����l�K����<孡��[�lE�T�l�������d�J�_�Ho�#I���At��W�����0��,T���{��s�kd ROt��b3m�Ԧ,c�G#W�Q3jҰ�}�ɮBC���ɻT@��&b��H}�s�M�(J':Y��tn�ߕ{T�D1��$x;{u���
��i�>�ݤb��������.#7z2���`8;\:�h�HG��e���Y'��֐�V�5v)�գo� ,M���	���u�o�)yb�
�~�kf��a1�8�����d�+A�H�\�GƆQ><�A�w}�=�J�<����������iN�M'�B�q���=$����\��s��Se;���'�
L��A��@��%�%57R�ߩ
�Q�8�n1EX�xɅ�Bt�w�}�F�m���1O@����z�/7ߚ]���#�7P�SU�Q�n{=7WE�1�iP����.=�4)~@���Z�[�^����lm̊��p/*͑�C]*'�6�{:`u��7�:���Pu�^�Ӝ�4e���h�)�������.W;x��
L��A���j�$ܕA*�j֑��w��]7�����3�#��R�1�s�b����w~%�l��YvE�ǲ��>�����0$Q���C��ΜP��Xϗ!�~�`׭�wY�,��70���A�"刻A�9���o��������`qN�����JH�] ��%�6�i_��_F�B�l�5�g�*�]� ��MW6J��J����-[ء�[�_��@�w���9���½�ぢ�����՗�s�����@�G�o{?=��D�y���˘owp~�U%k-Ia_���^=�h�Y�Ȇ�Y����
n ���V��O���U{�����t�P�D�׭�5�`EQCgK�w�${�I��į�
�ET�$|�}؃���IF��c�Q�"��Ip'�x�����xQIE�%��x�c��ݱF��`7}m���M�������?ac�,���9��:��Wڡn�qS����X�@r���/V%�u(XG�JX"�` �J4r��U��V�'N���faו�<����dK�DI�H[�����I�$f�u�:r�:�7j�{r��wBGC�)�(�g�M�k	���^�_x���zC��-���G~��]���
J�h��i=�d��f�	׊��"�d++���7���ާ\,n�*��uA��-�AAf��I��?��4��!���$�F ����w�����0��W�Mqd�yR�I2&O�XS�SO7�߿mNF:��6#t����!��j��2�<>���Sv�_��Q�Н4nМV���PXU�9l8ȱ]8nQ� ��c?L��k�2���"}������DvT�U�Q����wn1�y�S;������0�.<�hP�׍�/�������U�p�du����=�U���V]�c�̏�\�B,���^�T�U�t�X7]�R�f06�E��r�+�ǓHc��S�c�Ӳ� ����*�v��!��z�����NxyK������JF ��"���$��9bJ�o��9Sh���,��D�ꋣ�^�3H�g�F��Rd��"�D\������T����"_%]ݾ��Ҽ�.�\f�f�{gc(���>�r�d���'����PQ)7<ϑ�)���O�F� /�q)\���K���(\wq>�s���[�o�R~A�0"SN����n�p��g�/�n.�c�e�R�X�D��wtC�BB1��;��W�A^�3��+�����&�4	� �ڢ�e���kʼ�,5��œ���`�a�N�U��qQn���)��:>�N����_���w�6�1��z�."HJ�J�M����e'"����_Ӊ��Y	3G$zb��6�Ջ���lv�8:o���d|���B6�β(�t19�OOFr�{
~���IpR�O���N�R;��}�BY�-�V<A��`��ݏ��g.$�9z{�l0�g�}-c�u�W��.~$Ь��d_��.�m(/%�֛����O<WG'��g=���8���z��x^����Ϧ�\O��6���޼��59M#���3�ta�Wބr���h	�|��;��#<�n&�S8ܒ-TH-ǒ��k�	��u��m����p4�R�1�}���ü���5�_up����_�U�<�|�O��W�:� ��Rǯ���=����cw0�06��o���R���R��[Sl��IwX�u�}C+��v�*
蝲�*����Y�{[ٗ��q̲7^4���'K�B���o�W:�A����p`�E��9o�U`|p�M�Z$�Y��pa�B23nT�:�G]@���}i�?�p���.|o���=7� �u!0/���ˋ�<*��R���9�&9�U�{�#,K�5ʦ������x�q�y{�^Yx�V���S'�Ѡ`؃�-�/G:BDp����UWAz�^_D�8I,��H>Ɠ\ Van���e!t���j7��7��f�ݽ��(�������Ԩh�"�!� `l�y��r��5����|5�ٶ�=.i��R��*Kbb&I�^���c�А<E��@��[4���۩��Y�㥃��ae�G���_�������A��Y�[_i��yY��O��%tx����3�����Ckz��2ޭ�����M�/24,�8e�	��I2�/#��n��^.���T8&�R���ք���?*׏Y��ȸňHP�o��Y	�%�e>E:J+��E��t����[�x6��'��d�Rg��նV������o|�&�'CڝmM����+a|���i����aS/����Zl6�=Q��4�Lx��������;:�� ��" ���X�K��!�)��S�:���}n��M�8��dw8�D=ڹ�F��n��*F�����@Z2��Kc�"g�{�W���V�JrG��cl�,�I�2�B��&��4�4D�V��C�֝�=�AdL���Z��[NR�z3]_lӆ0!��*����1G��m������y��liRg�ߗ/��*�mt����^Ҋ0���\uDqg�{�uu{�k:���x�ϣNy
-!c�2�eR����?����.��{�nt���@�hڪ:y %E���/}\֏я�=�~���R��F�������D�b�J1~�fXC�7�2i�Z?���~=�C�$��r���!1Z�A�`���i+���uΫ��S�ed=8�똘O�j-2;�j] �[�?��k�?�Y�Jj��D� �s�IZ`1`1ɤ�?�k����Կ�h֘5��N��?���ꕡ�j|y� �qG�b��?nv��W�Ts0�:�$�?����#���$^�6H������#E=��n���ͭ�ϡI��n�=�fD�|QrI��Do#?���U���{{.v�C^q�
��&���h��l�_<����4�rg�c�Q�a}X��O�tчY�fmW�9n���K]��54��B��g���<%��(19�a���`��_.����]��5I�>���j����O������o��\�o����͙�ߐs�-B��jI�#��EY�ޔk�˻\��P?��$W�cy�v�����ۄ]-�5�*�
}����;[�x];�z����q���<��7ӌS�O�꧙�h��z�T 䍳r
;��.y��p����@��-�+����e�-�w�F��ʿ��*¤덍�ݷ���$��h\�T��U@�����?{=����g��Wtb������q�ڦ�A�����vi��@߾�d�㺙����V,@�*մL�؂�r��P��O�	�	����L�f������7чq�6���s7�,Z++x��e𗃜s�|I����8"�zD��T�^'�am������OT\��G ���E�\�qvAUL,��Py[L�;�Rf��oW=)�eK��4Ԧ��p����xC
>�\��+V3��]>�C��ZV�?����,=]E���a����w��%r�"�f���������C��{�t���a�*�}H�5�	E&�%p5+�yu4��u�k�yv�k,�5�����u"vƋ�2C�X�#�пDw������*!w7#��4���.~Ce�oT[�B;�υ�D%duwp�k���-t�q����ͤfśo�,�� ˤ#}�X�o������#�7�%+��Q��q�I��
�� ��2B����j<�-��H�m~X ���ٳ���!$P��i�`e���/����'�p�/vG]����oz��R��t����x�
huD%�_�G�Ṉ��l@���f�
���uہ05�l�?�����f �}��Q1�os)Ց�3*���2�W�!�����,����K�{�x�.r�>>���>����.��� �m��ڬ�w�R�T���?3dt������f]�wd���*��̺&��	~��n
�I�G>�/��^�yoQ=�5�����t�8d�	�g@�;��8����&�l2}�r!�lZ���}��_\�l"�X�аh��i�3>װZ�΄�Bþ��^1[ H� ���G�^���sb��PL�K��6Ǵ�<�N/�ܯ��p �6um�c޶oa-��7�eL�bH�{8!$���_Jc _����H5���a�a���Q�j�H&�c�����%(-6 �W����h�U(�:&H������FI8�M��C��*�ޟ��p2T�����ZvX祡}_�GR!��f�+�m+/��w̶� F_C��v&�����l2����p�O)SHPAO��}���ڧC�i_7�WT��z�>���[����2���Ep��^�x\��Fav1h5S��[��܆2�^�����6�.�W&��h'21D���S)��v( qȑxx:Z��"�Q��Ri�H}���z�1�����Ӂ�৞��tX�)s�/5;�Z\N�w�X<*;R-��F>f�|y���T��O��
�kEk8�!���ayIa��]��| �6~DS<Q�u��E�M&�d�Ă�U��V�pe�̖�|a҆�Ag&�=M����ɩ)~)L��F��K�t`�ܴA]u�m ��:��O�Bc
�2U�] ��^����/�b�=.����v4�A~���ovm��c�B�����ŉaI��?I��<��xy{i��J�F0�w0�1VU:H�c��N�7�A����#n^�ep��4R��v��{�
��9�����s��Td��W.u�8�Ϩ�FNI�`�'1k���	nt)��_1"!N��ks%�6�9�f���:	׈KD�q,��!��I�V!�>�2�\򪜭���.��m2������/M�U!U���������V�S���,��{�A�� 4��M���̓�"�6m��]3ᯗ����{���L��'�r�R��"���*�����r/O�s?��	`�m��=�P_����g�P��Q���8_�t,`A�C�{�V��T�y'��p�D���҆pre�}TT�f�i�\_���� �#^F ��S@JxϤX�^�B��b�Y3�q��� 6Z��v��f�T����#{�-��a?�LV'S��ҙSn6M�Y�ӟ7�'���&��vw����d�C������ rҪ�,�UQ�28�������ᶹ5=^j-���~]�sc��X�jJ�K�Y��i���T~k-B�-}JS��ѽ�
���Ɋu�)�����ˣ�>�~����z�g�h�Q0bG����a�}�	mYq��9���p;c@[ԓq�U��,#�TH1;�mdo�O�xKa�)�5,PϠ�`8�!��tՊ){�sX{c�8����d(��D�	���ȥ���驞�V��������=��<�|�6��=� %��rO6�t!�|<�f��|[|�{���d����1k8
�H�Ő��Z���)z��z8{�����J�=q�x��l��DDvS{�R�F��.4#�T��(�QA�Z�������[K��Q�5Oj��yYac�X���hZ�AH��v!�ﹿ���b����!�Y�ؿ.,5D�1�Xϐ��ϩ��wOw�=,�Ve�w.6y�o�F�|| B�4��.-�5o��ظ[�oe��ш�ZA��v���*�:5�]�B�U^�x�f�=�^&��X�Z�l��::ߧ��������~D$����w��Y@�A�d� �x��~��=R�R�U�(�p?-�ØV}R2����zY-��c���d(�s������l��I�xT��--�C�;�J(i������R�-�����L�jXEͺ�#w2���9x��5�Tʒ�����C�-mdx�	���ӎ��!�����C�t��yq�*�]q	+�[�֩���|'��f][��k.���:J/���?i����v�}�t �q4����]�5Ս����P+��_[�g��>��]�d�x���}.�E���kJ�?q��}��d�K��F���v)Ĕ���
 s�b�5.f/�r���"��9�l��wT,7/��ؕG��.t���q3���<�ר��r�ێ2ɛdk�g$ɥ+t}.¦�[ͨ%b:�+7rd�yb8T�e�<�J����OY4�@��V�;����<��Fz�@��ɐ��ƣ�~V��hە	*<-��f����hE.��*r��HP��h�3)���Ƚ�t��<f̆:�3�B�C�"+qE���tn�{*�ɗ�L�J�k2�o}��m�����6@�=ܯ�CG����ΰ�?��	_l��)���\A�җ;�	�P�b���>M <fT�����O�м�L̯OyIV	�u��U~����nn\��ÀD��N��4������*?�ǃ�>���U��E���"�d��!.e��}�i��p%J�����Å�z����Gv�M����L�?��!%-�8��v�FS��ʚ�����e���Zv�b3��^���ZP�+�6 ���qG�r�� $�Z�Jк�B������z$��&=��NL՘�,
�o���˰8%���I��n��`�+�ht��w�^z���8j�c�~J0�B8K�l���A������H|���T�Ю���4R1�N]J[�c¥i��fpje�^I�|�H������T ���hm��j���I��q�]n��a1@�m�,�]"�HjtC=�x���Ơ�VP��l=1��'^�v�S��;&l6�;�(�b����׌��1�z/W���b��8�$�M6����^|cT�����ۓ�*H��0�&8��J�r��X#�o�a��jWǸ��BKX@���R�+�?�Ռ��W�	�87D7�d�����х5h�N��ސ�m~RA�.��7!?����r3�����ї�v�W����|X��P0 ��7�컷������f��(�j���.{��B�	���oH�Bhf�0��kܘ�ϸ�6�-�u���ύ-���*ܦG3z�À7t2���\������Kb:�U��3zQZ��>z�Z���C�*/�˴�@Z!u⍓y���3�3�=nD�|���<4P5�y����w��Dn�_���wHc0)'x��&s���`aj��;i�ሞ��<yD�Zة��m���c�n��<���0��>"�,��v|3oU3����n��vd����	�����!_��X�!�=Ut&8p{��]�u�f	��ˬto�'l&-��f�7'�+����3Һb� ���dd萣!�-2���[S�Q
�w�H.���s��у��ھ�z��p�s ���dB�/��&���o�b$��~����QB-�I7�$��FKa��Ȝ� ��L�At��e����I��{�i=��$�UP�S�7j�﫫TGԠ�D���d�S(��M7�#��#�{W�L2�5�Q����-T.#߼�ț�*y��,��J��~����0�E����(�~�yO1��d��x�m8+W~�bhFP�g�Ww� @O��j?Wʌ��Wl
���l3�SN����#aUo7��T�TA�IA���/"�Tϱ�d�!�2Hv?���H���0\EU�p/��=�������NKp�<69Ͱ�~�Bz�����F����pm�hӌ�OS��ފ)�=���gZ�����^"�G�T�a�T~e�F@��h�:��d����Z�Y���q�P��y[��F�z����n߃�����nKR�f]���#N��?`s�((�C/��l:�T����}�H�����K@ʙ��a�N�NxPP���d)���k\��u�7/mE0�E����e766�
����羷`y�??F���L�� �"����̺�Ll���32�9��7��'�G��nj�<G��v����~|�?�ґ$��3��h�[���-�8��K�ڱ���.��!)��@nhG���|��8/�bX���OlRe���m��{ވ�����U!�J~5^�i�$���� ���l�@�A���e6dr���?�)��^�'/.��eTW<����1�]��{E��A�"�%�X���u{�w�����+U^��2��0;��6=�û��Ssk�_o���G�k<�T��3zqai�4�𧅱W��5�ޯL1������玌 |��,���M���v�П��c��>���UI��g����K�
_Q��Pj?�xdn��u�[����6�I�Ma=��6+��%-�]�%o�;��
8�`#ɑg4��{��nу?:�o� }@�Qu���>��\8X���\�OG~A�o����q[VlO%����I_p�g@�b�JMJ^L��!-�Жh�i5�G,�q�G?�t�,3�%����U��!J6��M��D^�X�x$��r5#V2��d���>Qp�{E,Y0��e��Uq�y�#J}D���XlxV65EB    f294    28b0�����Tb�7O����F�8;0'h
��i�^m۲�EQ���^���yܑ፟���Nu*i�GH��-SC�Y��98M��>�=�D\e�E/FM�g�v�~�C���_�T;�xA����:����k��ץ���l��ed���f%DX0�r�� �qR����/j�H��/�����b԰.�8��.ǴhVK��!��%,�.��֮oѿ�i�`#���0�O��:n��� �b^����Z��<��CE�o�	� ����x�D��ꏑz�7J?ly��uWz#�y���2Z����ۦ�@9)7��r�
�a]�7�[t�����z�!򪂭E��?H��{�1�6&:ː��ZBϿw9ύ�gӕ8������åt���eP߬��V�����"�������L�p/5H� {S�l�/<�t�5bJ}Q��^8M��
h2���X�Wg��W�sl������RХ�MN�p���^�W���f����^�����`�d>G6�$���~OT��	�q�>�J>�Q�"�rZ|b6=��	N�$&nS��E$���G�  c�yOم��@�n"v��'(���k��[O��������A�;�ڋ8��I�c�����]t�xj����1�agb���"�ۗ5��~0�,X4��sx?BZ�(���f�AF>z��j8�7pA[�����yi���h����(n���?3/4<u�����]Y�^�&����4��^�s�D3<T�4�X���c�i�{֐b[a^�b�Y8�{o�W,Yp��stnB�@�L�R_���k1 b�7�9b`��$��ܠst�Bo�d��x��e�������x/��%䣑1�_�@:��JQ��r����CB��H#���I�y�x�ۂ'������X���j�bJ��u�����c�_�ӁJx����$<�o ������]��v��9�����w�z��騬��$���( �Җָ�lia��(�����î1��}>��H�����t'��~�����iC8x�j��e�ZQ�����,�6h��o6��6�7
k�)po���Q�6���'�Q����%EL�tjշP!=p�D�]w��OUr�~f=��:�u��k)����5ܨċ
��n1ȪdB�i��`6n�����H~�����h,; X�/q�H<�� ��aD��圎��e��r�'%g���o�`�/"6�v�x��w���!�do3����B�|�F�D��ٲ,	�y(���w�@�dT|�����D9��y�H��x2�V��Aq^��0�Ɨ���W�w'o42����Ƃ1�����6�DQp<��kF�Ͻ�uԤ�5�V�{&XϤ�k��4 �� jr�W��P#zɥ.���r!w�xEmą��a? eĻX��+�'�=�Զ�-�X�)	>6�����R0�Tʨ�0�SI��;�5���8�p��בs�<ǈ�F�c�om :��)�HIx��wI��gA8KG�*l>�z��L<�K��5#�����&xe,(��+�N`�ѱmoP����Ò�W)а�� '
�&�%a��0摐�y�M�H-��W���pk(Jl�	D����[\�:y�������/_&!����/iF�5	���nZ�F	4 "�Bk-ۉ����JR<�[��{@��csg�2Lj<Wr��Β��7��~��I$�b��j~K�wk�òh�2-'��f��\�[�Y�i����$�:&�^�Ɲ�^�>�_��B;���R��Ďܫ-~D�k����jwi����q�����b(�������~A�X�b1)_��aC������YT�'��vs�1�0F�*jߖ>zI�R�7����������s�ꅓ��#��$N���
k������r2:��I�M�0�>��n�#�2�'H�q��9䐵���p9o��^� ��%��`!��t]YZ�-�52����6�4��sֻ9N�_���#���Q'�N�����J����O��˭��W�sX��L������J�FD����z:fP������jC�~c��M�	��#�1�Oַ�u�K���+��Z	I�f�?�0�'ߤ��UI�W�F��������X�(�i^�\�]J��RZ�ޮB*Tl�#������`I�Q���ˮv,@t��������P���9������<õr�q!j�@��=WK�'H���Ā8i�����Ql]�)l��K��k���́�e�ϧ@1�bBk�
�`ڦ����@2�����ϩ��f�ȭ<EWX�<"�(�<sB���g(���Ⳬ`������~v�?e�Ƴ��}(��ZCVà=O�U05�_����ص�dr:�qPHƓbVb΀v�><N:���(I�%x���3�*Y�w�����(��"X;h�B���8�߁�����j6����!��r����p����B�}��[����d#mN������LJn@�pv r�r��,��w��gB��@�d��>��d� ��i%��e!�ŀU��jU�q�J>:I}H_��񲸭\뉴��<oÀdZ];�{��f�]$aMp��&N(������壤���VAh��i�`��0�<�vET�Xj�[C�S$���el���K�N �iș����)��uΣ¸?z��ﻓ���H���X{Vl�K���=z��l�;�HN5�!���^�=�h�DD��=��f�N�+y��;I�j�<?7��/ѼwZ����b�Go�IOo��(�M֑{����n��䖞(��؊����l�
b��ʝ̐W�*U=�4��	�RH���È5x�Y�G��0PD��V����eY�����s@>��"���E��e�:��x��`i_w��c"��F�26&�A{��N,������0�eⶹ���A��f�%�����u�� ���l�������!b����U��e�ճ��]�V.�7,��3���u�ˤ`�z�<�
F��ٖ%�;@��C�׺�^�k (�,��O7,|Ƶ6��l�*Z�UG����-�i,u8�_�nؿ�ֿ� � �u%T���^~��Y����8���}���Ez�ǝcoV��,�(����-���n?�.!=��loF�_Z,ʛ�uz����|�"�݂}�'�֜�TZi|_�	�Cf��"PP���;i צJ��
�Bp��M�fI���$�I�-S7�۲��}a�`�LT��č���&�k���
3)n>�媶a�����*�`�|�F;�8z:���U���7��'�_����c���,Lj?��w��/΀@�����Q�O�A��ȧ��g�z������6z&��(/˩YiI�,\qφ#�h�7��2B��{qGX΋4��3`!C��d���**��g�!�4M>ET?���_���@��ϊL1�0@�[�˴��vA�������peT���S�(DH]�47(u=^��~��Umej��.x�B{�l�֜+b�
q �,��I��b�Y3����P��j�z*���W�X��(��oՖ�M�Y��g6��
�Q��J �3��ܲ}cC�BЏ*��e�Vo
���P $P3�5�E=���	��Gp�c���3���})�����.�{ʗ�`��%9m�"�^R��G��3��o]':�'iQ�yb]v�_��Xu������rC8FR��+��\FǇ� �	U2
�"���B����~Xb����ZGJ1Xz��1n4Ȟ�1��1������ږ�Hc6��Ri���H�"F���;�� ��Wq	�W��Q��Q��B���������H
�S*�tI;
�$��ۣ�x��vs
�KC�5�m��L������SP�-��Px��t		A@6�l ��gz�f<���XxLu�s�m�&�X�m���25���$��p�ҫ?b�!ԗ���+eD���odT���a���c�6�7�r�8���[�Y�7h֦U�Z5�ț��S���TL��UP'����|B٧��}�f2�nN���yJ6� ZpOk-��U�(��ֳτP�;�	T�MJ�-��5���(�Ͱ�����&����*���S>hs���
 (6�������2�y5�[A#�_�݁���^@I�&@���3����:�YJ�ێp Iv�6=��_}]zD����GP���Xo?D2�6,_��N'>02<��
Y�D��$�X�'��+k�l�s�ټ�s�;m��E�x�1�0ڨf����6���Sb)?+ �oϦ�
8�gF�q���,/E* �P�H�@��L��{8������G^G�����Q�t@��]�}pxF&���)D\� ��`���^cy��\�뽊5�u-��{�\�[@�F���Z���^3'F*{{�q�y����H�܌ܝ�m	��p�;��e��j@�P�f$ZY�n*^���Q �� ��R!�w�����Ű���8G���Nhk>�0/��S:��)�D�g?l�D�����*���Py�\iL�[1��5�1;�����="�]dOUQ��t�ͳ��t��u6�p�}�e��&�QM\L[V��-�Cg~���� �p}e�Y6a�F���}v�9�Jm�A�n�0� {�'@G(�P
 �a�~���f�*��~*I���tX��(�T	Z@�����	{*M*A�,��j���x�8��H/�e��:oޓ��,\e�w��B	�/�J�����U�SP�ђ�[1���c�+O�= ���{14O�:w7�����B�, �D1� S�d�%�my�QJ���I��g�1Y�� �lu�/�ܥF|�J�,<Y�/W �V�ߎ�\�"��(���v���@E�HX8�
�R�mh���2� =�b��Ҽ�K��8�C|�?{3ăڠ'J=��$v��5k��`��/�n-��3s�iv��F��Q�&u*���O>���K��v	�"���Q�
� d���!�A�#ĝH��D�DvBZ����2�7pc��RFٍ����p�tU��������d���?�s4�1�^U5	��@�z}7@�2���.��>�~
Ǉ7@���5u���$ʟ���b�=�-V�@0�H��.`�)�g���/�O�&spF6W��S�LP8�nJ���'���ɦ��h賙��JD�@V�:\�s#�+���������#{AՈA���^�ZU�(��e�l�w$�5�d� ��p�FP��!}KF�<���y�BM�h+�}�u�C���k%0�t�
�����Ox�t��}�G��52��)��m�#��=�%$WՀ��2�q���^&
RӸ��`v9���z�c^M֎�;K�D��7#��f�F���:�a�{�<���<�������B`�|(�,�Z�~-�_�	�H���M
�i,����;��t�5Aϐ'�7[T{�j���l�Y���Ch`T����<p��qE��M�}�):_cЇ0IXD##�^�wu|�̤h�1Cr��qADM��8����3��;�b��f�o��	޵��"bC��\�`B�J��}����1*��	ry��fF����1o�a��!��ˠK(z�ӽ����"W�^����JTj����iu�㤏�+�~�_6���+�LY����59�ϣއyS!��� H�:�\x����a	n	-T���yI���w�:��2"���T��.����������q�0R3�T�P�m�UѴ43.٫<�m� t3���AC!��g�_���=��8C�c	*�6V�;�T�LZ�g@>��Vc=�x
��c�Svt"4FT ����z�vֈ#+��\�CZ6�$s,[t����u���=$�~P��i�|��>r�&H�����o
6+$.����;�4x�z��gn�*�mc��m�L[�d����H�/"��$��y��i9�?v�zV�F% �q�%&�ʣ�m:_X���s�<,�*����m��J}囎�0�H�	�b"���յ��H��9�h�oE��z��Wv����G���6�[�AG�NyB���ii�&��������?��S�K�b��6�+�ct���@'潜����]�J���Y��cK�Ԥ��'�%B��j�V�T�&���ji�&s ��K��d	 �@���\���m���������foP��NLM�p!Li%�B|]��\���z�-�{>6yʹ�QyoF�:�3X�U`�3p�J��
�e@��sݝ1øڇ�]���:;8������Pܭ�J��J���1Ye���{ڿ�e�z�ҝ*�հ:���LX-��b�㯈��B�c*��-���"���_�[���gW��fEtU�k��x��W#���bz⢘����ӗ��0@=ǘ�L��竀���#n[��ۈ�'�������:�pB���~��ǫ�ㅄ�ɢ#��������Lр�A�2({��L���A�N\�ZV���	c�%!3����K�c�B�7�����9���	΍��'�M����;ΡfPh�e���k�%%(���$t�������5R6.��_��|t�g�}ְ�:�J����m���4=<��N%�.ñ����3��[�K�!�ްqO��O	>��/
G�-�EK�"y|� �C�&b����3�t[X�X���4�o�2��}l��=4�]a�?��.��u��F��;"�9�L�����if�g����Z�3�P���<�.-:�>+�?��gt�B�m�ֈ�i�q&���g�����d,�N�v�0-*�7�ʂN-�'�#��m x��/��NF1��ұ�
������G��ê�nD�{*�-���
����!�'�+c������QI͂o�Y�T>������>God*�ݝe4��1p���O=�ʕp2��L�QT�̂5J�� Aa��������3@�5�س^���h+�_�����no�e�\q�H?`�ɟ���X��4��¾V�&$T�?�=���p՚�#T����F�-���]U��޳)�Q
����F�gH�T&�Qk��j%�cW�� !�'���r�_��_�ll����Q���[�x`N��*������2�G������p�W�#)�0�L�`6%����.4�]������>Vrh>���d�]�<�q�b ��q���g��g��[k�y�[��/E�*EI�6N���23���l��R�O��^�"��TY��B�n 7��\�WN��펈�m��!�9�%𴹱{ �q���0���_�~���7`����W��i�{A�1\��$!�Ɗ����(���b�M6Kt��ck�Fݟ@���Df�=�_��d�w5���κ���b�ì��Oܡ*� X@R��F's5�6Az�{�q���KB��� ���0x���^����__����R|�k��ֿ�-���m�^Pg��$��FZ���m��z� Kٱ�.���)7;ɡuq�3�R�o������Ʀ�>������t�b�a ��G�o�����D�%���l%"*6��:��I}(+���3�4H���\8wR�����S��
�K���V�E��\(R-�)r������.;3��]�-�S+y\t�%�M��B��%������F�$���N~:�s�nSD?����&�lnh�R{u]+��ǚe�]�g%$"�|�{���[��U�80���|՘�3P݇�5@����!J��S�óS���߿�r�
�9|t�������:�v?]
]#��Z�<��P��1���9�~��)�O^�]R�:,=��K�v��۽�|�:�J����'N�8�|��&�?��`"�J4�̙���D8FG��|PU�d=�L�ns�7��F|w�o{�W�en���w���y/c+8�C14������Xˮ��PJ�|$0���kئ�@�S��3m��Oܙ�H�7x�[�8�l;�l�*l��'-#筁q�NB@�gB�j��e�'bߓq��ά�f�!�	13iH,��"A�S�#:d��;G��(������A�zc�8�_�Ƅ��%ŞD�"-���$"�$=�n^�ؘBo��#"v]*!c#�G3��]�/V��qNE��N��`ao�8�!�3S��H�H�%�b9�s��
��5u�k
�C?1�?���y(���|EC�M$^?��F��(�(�̱a����9iQ�?X�0���Ҥ�'�\֮RgqN;�dH4P�;��vZ��܌I��p�"�������~�I
�LܘQ�K��n��#�p�jR6C�"��(D���=_����-�Ƞ��~� �ɖ(�SR��UE.�;=fz�}_�t'	�#&�<����2@�-�ʍ���o�@i��L�Y0���
3�E��e}���\α��.�7/�� �7ۉjȗz��(�mB�ٲ.~��R�9��x���kL�N��Z�������9r�P�'E��Nq'��J�E�MOӗ��
�>���2���Y4�B�N �[X��0Ʉ�?��cO��P�)�����T���΍ʱNo�\p5p�����V��*Y7G�<3��I#vۑOd���a5���rh�UV��A�?�38��Al�Fb�P���q �ښc�j*����0Ѿ�|t_o�׹�"a=L���vz�ė�r�75
������"�;�4�a�L�]�������fi�\�FBΌ��]��c<|
�E�w�g~y`ot�Q��]���C����������B3�o���9L A���#�*�1Pȧ���m]�~��{��"�vi�Y_����Q�qFÚ��t�~������i�xu+��㽓�=8wh�l�f���`ֆH�8��G�쌚�F����)�P�0ǒ��6�.5t>!��H���Dg2�-�p�@{�J�CǉS}�[kP˙�Q�Z%	[�xxS���4]���k�茩�d�vIr8Ҷ�?�i.�^H�Tp"�g$C���^�`)�@�u0���{�~�s������<F�;�aSd������~��=4Ud%�����i��2W³��b9��k�TQ����j\���ή���]x�?���U>2�SDu�N���O�������6�MS��yi��@x��i�L!l��;�H�O)�V!\��DE~���k ]�uV�}"� �5gQ�\�B��k��j�cd�.zr��T/��e� p(�!�窿����2�Z��n!���6��&�9}q�m$������#!�%��ye�t�� �c��1�ւ��-k_�a�X��>�n�T�a�!&�Q3&�$ȼp�2<?\�b'���n-����d�k䶽V�����
�:�lI��2B̈O��&��m`h�[!s���8�!������-%JxB���˧��:�����,��fGr�6:�"uEVv����QKn��U�64ي�C69�3ݺ/]���j8m�/y��'����JHn�*�j	yR�>�i�w�{lh&��������� �����j��M��� .�`JBo��(]!.��H3����z����kT�^$�H����ʑsE�\����E3��>,�)"�]��h#�QF����(Ş
~��@m�Q�#i�������@NS�!�t��d�.���%��AL�N�b&���WL߉?�	p>g�J5�}'��@w�#�T�r'�_�6��(�6���J̮�|�S�˶��9��*gk�<��F];me�҆ߛ1���e@։G�Ш�L�t0oo�5�A�`{���V�e�|Y��vrн�4��oc�kwn͵`�� ��}���9↫���a1k�+� ���UV���	�(�04A�c�S�C��'�����㏼�b����vw��?�'�>�����y2�<�+>�*���׏��L����ukr����vg��3^n�j��/��}�h}�L^	8�Yf���ڱ*�6CܐAg�!B�lwۆ���Y���}3uD��)�S�̳����������������wk�@�� ��C`}���|��Vj{�t�9�ğ���7l��;�
4�@e
Y��	ob��Cs��iO!�ݥ�h�Ed�e����f>�z��D��1�S<@߆�CC6��u��⦔y��T� [黄 ,���eK쩲�$U���9�{�)�;L��s�ֹ!��L��}%��-χ�V�<���
�3�Gv`�Nsk�?!�6ן@a$xf��1��y�%�Ho�l�J��F�V��9,yD�Uoڽ%�'PU�AB��j����4?ݫ��~#�1��������`�f<��l�t��!�|�te���B���n�̵��_o��O9��I�ow�C^Lr|n�R�B
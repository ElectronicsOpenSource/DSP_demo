XlxV65EB    fa00    2e10G��������8�u/�YZ��p�	 ����l�����&K!�؏%"x�eP�n���Lr��ncX�qF�]��^j0�=n���tY�>-�*AM�k��6t����x�ʌ:`I�j���b?��t������������*�C�Qe�ϯ�7�i�&ť��5���jb>��wO$���1�@��5Vi������U���^|b��&�c��aK���<���;<'dOg��kE����B�u��n�y�-v�p�hk��G��G���9�����w"�}ĸ��*��O�[U�L"����Ga�P
�z��hm��p���!�IQ�6�p�q�B�}�4�n"�7��[>֗�c}7����0�8<F��)A5�����G��r��]��pJ$ Z�C�x�i�C����W:m�(B����y���]8�S]v���E=@5l��3�@|�h����\��	 qs����8v�l�U�#�D5%ܿ�Kt����f����Տ���ک��uA��764~��"I'���T��)�L+���2S�zCS}6�}΀�W3G�(�g�l�n�-�Я�8�γ~���P��Ǌ��ʥ�euh�?i�58Ȫ��s#�ve_7�D�	��(9�up�DE�;2kB#Ps�ϑo�lB�B��ژ��GM�B@9�T|D��Ǽ�a��q�N���f[�H��jO�3�T���҉�>M�"J�'��X6�M "pj�:������-������;��-y́2���}1T��t���L9�����w��B$d���}��BK�JOs�.:"O�^�GY�'�&O%�
6�Fg�jF�v�����0e�ŋ��;���gǯ���:uZ�⻝�L��$G8N���/�V81$��^�2����� �V��"�1{���� F;�yH���xp��wN�(��{�?g4�ɝ��Y�@��p��*s壼�
��7I��3��u���`�����CQ/�.�o���v���c���χ�����-ㅂ�ӫ��jN��@�ܐ7O���$��3bL���=^���>�?��.Dy�nʜ�o���+�{����pk�����b�����vף�X |6�D�'[JB���Ħ�V�Ȑ�t�Jm]��>G�Iķ���m�ߺ��^��h�f1C~Y7�# �1*Ƀ�_9X���/�*l���h:���幱 �f�qx������7R��L��7�70���׹�'Q��I
��֯a�����̙,�����#?�Ǆ��,pA�A�����We��K��A,�j}3Z��jҔPZ�t��3+]u(�tJAd�wH>{�2�H��g_U���Xl���R��To���xF-����(Qh��J��ml�W�������#��6�@�?'��$�0֋����ԕ�8��+i��p#
��	��ǥ~K��F�g�kN������R�0��Q����}�/���5�?��!�VP���&�6��4S�k�*�z�N�A_���G
m��P�mvn��c1��΀�%�ўc���3w�(� �R��EҢ∬�wH�����yG �mV�]w�!#�w	�5���*�ɏ��|g��{�t=���Tp�DI�s0�^��9Sn���j��A_�pА9T��!�b&r��\G��bFCA�^�LINr�+0Ց��d����&Kꈊ�B�q�14lQ��N\Z�����O'�,�\-��}ڨ���|���{q�`��{��8����\��Xn(վ}
E��T�a�rRg��i���Tr"|L� ����k��~$� ��T9l���9���%&R]ÅUf��K��Nr�gW��.������GI���D:��CfCF�9L��Cd����Qh`�E9W��M�����{�S�7E�X��� ���g�*�)5�NQ����u��͵9i�2�Q���y�Hkvd�J���(�z�04�B��C�|��i��Ӻ&�~rf|�G��\*��H�{,�eg���L��n��s��P/�ƛ����s���Es#2,�؅F���E��^_�/܎�X$E5K�S��S'cG7�	�c������(1���!�t]j"�b����2����?:��4��am��l��@-�A���畱d�$��ۡܡR:��������F'��-4��R�T����g"\6Ǜ0%s�����'��J�q���7L�O�s��oV��u,9�z�(���f�����u1f��<�Mo��b�a1�>��wj�!k�2�5�����ݶ�\*������h��l�t�����@����na�;�`��B㞎8 F����!tX�>;�����ܩ��86�>��~!؅�q���q!���t�2+�_9��u�彇W��n����dˮdf]!�㌇�KUtf�.�ΜsA���������rDG�e������n���6@F,�C1�2C��/ުds���&�B�im/ģ�yi���p��f��Fmd 1�31kO��W�!3������A�eA	
��B��@,�g���]M��_<���5K�U�K�[Z������ֿ�UK��FuA��*��m�,msF�e�]6�x�}��qI�C�J��d�(�t?%q����H%����n�vA�/e7'�V�R�Nّ��w��G��Y����#��H�d��fIj���Θ�_�$R������i�����с�k^�c���ɍ7I��q�	M�I~@hP��6���s��SN�B=�j+�C<�
�Q|Ya�]���mJF�%yP����7tNa��8ٌ)�Y�Ҽ9�Z~�oiA��������B�]Q�e�����i�������9������*�.��^�WZ/��,���9:�2���sY�=v˃"g@tHRj�y$ � ��?�K/�#��#:�ב�;�w��k� dΘC�j� m>M"H��bJ���p(01�BZ(#�w�w���%?�C�u�d� ��ܻ�ާ��B�b�J S
��qZD�f�o���H�n��e$���gێ�ԪF��0��뗑%@�UH�Q��/���r�g0v��w ���j��o�FH�rU��M�h�`�϶�M�\��w��T�D�n�$Ӕc#�Qè�Gc����MjN�Qz���d0��B����F'���^G�֗�"3��ml���|K��^Zn8��$��cRB_�N`U�-6_��Vf�5� �S�B���Y��S����b�fN��Zd���<�*��1�bi/�.#:���>��e�����+�]/�������	�a��ۜk�!�u�=fi��s��F��Z*V�~^J�9�~����(BX�	Eg�8V`2/�3d�`�;v������(�c��a��ٷ	��-V�����n�4�y�3ܢ�.��`c߬�ե~��)0�ώ <�g��q���7�n�cU�Kl3�7�}���@�jJp쥀��S��ژ���?BJ�F����]d�HW3?!�������.�G�!7^�і&.���vrop�J��6a��K�T�-p~��ȱ�̭�`o7q�����f��$l�����pg�<�����F���'�w�E�f�;����͂y{��p{բ"�R�zMR9�K�ܪ �C�7�D3H�XM4�����7IN�c
'�����r�Z�}JN}0�{�i�m�u�����p[O� ���H��s��(��9�a�K��G�k��?e
?.�D#x^�Ҥp�aE��JK"�A� f�,6�E�L'{lZ$�ts��`b��ȹ�o���A�0�\Ϯ�9�+�C�6��b�y+�U#�~{࿧-�S�gڶH�5P�d�Ik��P�/���:ŉ;[���E@Orô�!&��,�D�n�ݹ��$]�y�	�D{Y@�5ƼL�h�j@���5����u��UC~,�O_���~G�W+"Fs�:e�呤�]9�4Ě�O�n��l�)�c ��S����t�l�.ď�aZህ�۶�	���TWFҡ��P?s���r�.�r�B+8�	�:�)�X��r��6�j�x.4i�kv�O6�}Ao ���5��Y�"�fq��'P{�������E6��t��D�k�t�OrD$LB��$����]o �L���l�viN"v���� �p/R��P�8��Q�9Ц�W%M���CboB�W��8�n8L��M~���W.T���'�5�����&����N�Z^⦧[��&+�c
�.8�>�r��o70^�7�Rǈorр�qi�vgӼ䫰7DM��8�>>6����8	��A�/��;ϕ������v �ޫ�P���^.|F��!$/}����f���L���W9�,���r���+�)2�����G��.��|��I���H�P|��Ԧ��놼=b�ۿ��">���)2.��������#M��Np3뛔V�T��k>��<y��Z����W�B�˷o!�(�L�9���>��U��idr+�RA�~�"$]CA���*3�I�1� 앑wE{VX�Y�h����������m��u�k6I .-���3�)���~������y�x�|�.�������n���������0�K}({,�O<�}�&`�O��(2� [k�e�?�ܱ�3z�z*���Ю��٪�yf'������ #����L@~�0!�*���a2�͎��g^�+Cq@q�吻�Ì=�Qk���*�=�fN�\�xvyF�Ii��K5'��(��!N�S~����]�g�[Y*D䛡ہq��3�臅��9�6<��,f�O�I��4/3�_Of=��EA�d!-@�^�a*�L}�i;��3�%�n�W=��{��M'-$�:{�R���%��2v2�t�k0��l�X7�ucD�#�"`�{�)m뵸#(�7q��)�� h��C&N���&`����Y:>�z�n���ݵ�yp�F��q`�}�:��;�*+QW�K���
�0��	��ePq�H }X,	�Q�� ����%�$�*˫~��y'�2!:�Emi7�N��l��\�4���;��-T";�,�i��^����/��WRm�����Ƅ!���FE=!p� Heg�'���̄I@ 9,ƆN��c_�^�}#��Np�g�FXNYG_�e��圕�2�o� Xi}��jC�cv��氿��Y�}g&�д�������4!{7�k/�[�`Z��ː�����^l.���ҹfjL#�S/�|��͑ļA!��E�m�@,�s��&�ʹ��H�:|�?S�~��M0�P�`��%�#�ϯ���#����	��~�f��Cd�H����W����f�u�ڞoΪ��'g�%z�Pg��|�L�ą�a��k�5���N�Q��bG�]�dǮ3������:Y�<�Y�,�Ŀ�v���I��nH��vU'N@�Fw��Dk|&!&ߣU�Ò١`���2���:����A�1u�]����'�~��:)���$�BZ8�aI+J�2��f��/���ךܿ���o�1<|�ɸ6�T�]C��/o�#I���
YMs��B$�̓�Du���@P_F	����v>a������a
�;#cؙwZr��<�bM A���(
���f̍� ��}�MlH�#�6 8���E�􋒖aQ�����v󀐛�L$�'�w��z�������r��~���&���pVy�T�l��{�cޭf��:��Q쳿c}=�ø���Pȋ.U	%��c��e�sZ+�����+-m3ro�0�؋u/�,Nq��)���A�!`�j����	�."��"視��`�?���>k���:��sҋ�*���=��^�_����&�U(I$�&��H[]����M�XP�vր�k�A����8#jC�p*Ҷ��bh&�U,��)�R�Ir	��bN������e�G���U�Aæ��1䀵��)������83IϷ(�=h���	���LQ������= ��.[���nLm�<��-�woCr�|OH *Λ���`��,×��'��C���`��C/g�O}�c!K���:k��e�YQG:�Z���8˖)���|�|*�CጡT�G�}�k����7����鈤��J��E��W�2A�I��п��H���;D�\�<�f�i��X�v�k��,)��-�F��a0)&d#2z�W1FY�������Yzj~��J��=G�`F�M-b=��ãv)d�Yo�h��⚲:�y(�a�E戌���1k��!s�:N��M�<�j�+3c�᯾��V�_V��b��XnT��	����Lq�w���!�������΍���$��J �Ec�\z@H�$�82F�����:���Mq�-�E�`�������7�T9��0b�7�~i�!�,���1�9ϧ%D1�+&���ttrN�nX���}B���]��Q��<9çM93Rw<a��4����#��g@�d�1�ja�-JF��sU��.�@�,����N]�-��)�Y����!�Rd�!����!�E���T��Iۥ�Na̪~�:fbJ�:N����r9�0B+&�\4�.g
�w<��`>���kl:����0:����3mFhq�VUL�ZNn�tk� ��x�!M�(�~����84�HiO�����r��O^'��.zb��2?J�;��P���"�O�构ݝ[���x~s67�ґ�Pר]F��3�h�ϩ��
�<��<X�-�c���8g�Ȥ�����|�����]�?'�1�5��T=&d��������>�_u(s�k�7u�� 0�1d��<(�F��	�t9�OU���BO�u8%�Ĳ-ϡ����ﭞ��M�2�v;;X��bY�<�8�		�������o�=�����-�׳�4���|�[��7��ܸmʸoAl.��}DHq0xC�Q�|9���Z�1��IeS����1%�P� ���6N��Q���Q�dG�62��H�vd���#�FV�.~�9�`��l�B�D�7��%!���Wh��	u I:+`�|�Dh؛��{�E�����R�_�WrI��뀃���kC%�P;n%vK�Y5����C�+�\�����l�6M�\ZT��8���_Z���S*�/�)K�B�e��mC>��D�.��.V�j��C���K���Z8���FO�X>kd%��7"۟
Z��r��(�1ԫL9�{N��#��\�sã҃��"�ƛ���b����")�N�����h�z�&1e��㥺��у@+X�hхt�1�h���ځZ<1�$PjX���n;�K��J�{��>XDn����M��q�8�o�F��g��l���[��ԛ���T�,��G"�ؙ#R����|��p,�g�Nf�o&6УE<7l��e�(|���}�/�	�@"�~-yPp"a�d�\�D�vJ��������h2fQ�)&��M����R��ŨL/��QK\CG�_�£�c%��n�s�fO�R�2ˑ ������:���s��Z��CP�E�&���B��R������Od��Kd9���J��=!!G�y�O�#s!~@|.s�J���#�e���)�ր�;"�m`9+�]��Ț��!݅ႆ�2<��r<�t~�e��ad��fq&�֌gܟ���2N����"tّ��D0�?2�0�lT�|�5���sFC�.��S�VM��̿\,���ъ�ׅ�դ)|�Y�+1Y�c7� ����~cam�%�3�?x�^���,c6�x?t�0�sAC������&�B�}r�%I J.�����F��W$�Ep����.����XE�_4������b��xh�]\"R�T
k��-"S�5,���[�t-��pH��Gaq�0��b�F����N��|d?�,����9�&t�CSl�Ǝ9����ғ�)�15�FMsm�\CQ�]�?����2d���!��1���fw_}�����r<8zY�0�������0���I6�s���=tx0]D�ۋxD�3��P،���R'ڊ���E�U�� :]�d@�z��2���q��a���n�@	��k��!M���R���_���؈�;��_UAL�K����H���+R�δ]��]uBB1]6�����wT���s�ᾓMg��i���M�8��E��R��q΅��f��M/����.`��we���8��+�����¤RK���R�'݃Fp�3ɩ��y#�39�K�{�\Hl�Y������IB�A�^�w�Ua�j�:� ���Mm�\���<�{Su�YMj��*��P���v���v����댋P�%�#��!d�i:Z~&2�`|F�Lk�S���<#+`���kr�� ��S5Z�����@8�^%AT=J����h���~��W�~"�����j����D@�жvq�E�(RUCȜ���i=2p��5 Zj�����q��4�0.���`��/
�(�¾I�,Q�;�w�]`��vhƹ�*CB5�=xur��K���R�1�CX����͙�RlZ4�r��,45�3b��H*b,���#�-��҉�#\E��i����|+�Z0��3X�2H^����*6�E��4e[�����y��U4��~A1\�;��6�� )�J��(�� �)��j���[�I)u���%�1v*�F��b>KQ����O K��N ),ʴ�x�����wq��:�D��ۼ�����t�ƀ$V�H��'Bx�@;o\evnϿ��a'7pv�a�L�W,�p����8fg-��T�S��&�Q���In|���We<�v>�Un/����w������zX@��	�����&��u�hN�=v�Ŀ�̲��F�`Wп�{ObW� h��t?����׎�	�����J��RK�©�d�1d99Jn6����˴����u�?Ab����8S��(�3OT:7ˋ��+gݪ�Y����D7���1�/�h]*�,��BH�&|�!�$����`Bu�k��<�|�2��Q](�i�Km�F쒳��5�%H�?{9#���	� I}@y������
����q*����e������WJV�g���kI�'/e�0��1��C���_�5%b0fn>g"Jch�Ц�O+~T�	��aύ�i8�_�N�i*��~�y�5)ǋ��J�S�X�����.}X  h�|�H��󣠳@E��-��G�%4]���O3�	�n}�A�ʵ��LӗM����d�[5)}��jU�����F+����獒��FWע��Y��t@u���1��aJկ��.u�n�)����	�Z�'^E~5��t�aO�-k�eڝ\[�[��dRVb0��ns�����q4�rV�KY�'y��L*��4���t��_ݐ ��,b�G4y�P��W��h잓%� �&vg>����d���M������Xz��y*�26��΍+= yGDP���h,;�Z]�~Wb��S4-iWY<xҢ�ȶ�<AC���Urߠ`f*;i��R���e ���F1I�Qnne�<l
���V���M���7�
����ڂ�D��-��Kq��)=��fT
u�6��-��+dl~m��spT^������n1�w׃��ɘ.�5zN�Hܫz�OD��yl��M�TM�ڸ>bxp(�)|�#� L��n2讋a�����p�d��y<���x�ͬ�)�t����=� t����2j�\hKI�\���_;CF1ze<Lt���d��*G�
P.�r:N��w%e�C���W����l��D����?�*��ф���b�e��vR�6&����^muMw���C�6t*�b'{��SC�yV�w�#u���J��B�:��$&Śd�	�}����`ٓ�j~(ad��%Ъȋ���c��%�V�f��ۄ
��De����]*Z�^SmZn�-ܚ"��!{�^Hy�"�&���-ޱH-�f�R�ÉRp����S�Gx�MS��}S��D��2LS+��p��r��o�M$�����M�O�7�$H��m�U���Z`mx>�ۛ*����u�d���K\q
�)J$I旕
��Ҷ
������#�W�E������C��&_t��?��_�L�яH��CYE*0./��9Ie�fʥ��f~~���Y<��bSw�� ����CG��k_�����),3<�a6 �S�h����ZuY$�͚Hߗ� $�]���U)L$�X3�V���X�(ĭx�W�V5��y�%]�����vӵ��Y�aE7	|7���b9����n�e�;��fR�:ĭ���-h_��>8M��R# �T�q��\v�o$1:���^�o۴'��z-�xZ]B�H	 {[�:�9�����*��ԭv,[��}iì	�N�{��幸q��I�q1��u���6�t�6�����Kc��3��v.�S������>msׅL�����\��*�'��z!���\����j�6?�{�7����U���ql|�q��c�J�&�!�N[�gi]�����
x��W0�fQg&h���0�5�G�w�֒*CC�p} �f�� ���yW��a�4��c,�Fk:�S��>��#�8����3��~�����08aGqM�S~_t��x]bl�98��g(�))C����6�m��%���ԙ�vSe���&K�!v��g}J�j4����jW�;]����f=[oWp<f�SK�����9kb��wCs�iбj>~�Ww�㮘�R�52�Mo9�b����k�5}�O�+�`��O��1�Mᚾ�N߂��E��Ц,F�@��
c4`���c��,$�ƻ��^�e�
���;y?�Z�ċ�j2���8�2�g���/�p��}J�We�G���=S������h�*;��h�0��=ͬE�xQ�Q�eV�I�(�5b�ׅ��$���Y����4�����w��0/J��e1��Yi����������`6���<�3�#l���	����,�/�29�˯�h@��y�U�����rF����縣�ž��	���m��B���E������m��{�S����P�R��kA���B9~��̟��P;n�������(N�z�Z��OY�V�	��>�g�B�9@�$�
z�}�*e�j��YR��"(3i"_�i�4zxe}a+a�C�P�U�Nf~�����:A9v��Fj�#C�K[IU-]�+��L��(������y�,)3S�Q���d`D3����H����c�\��>PP��Dq�!��xe�5���������_�f�]�����w��s~�7�@�:�?��T�������,[�9n��������g�8�{��`��.�B��e�L���=�T��EQJb#3�qH##5�ʊjQ�#�$��}C���h?��>S�'����r��,�V���o�gbt��J��^��3E���l�ݸTq݄6#�u�>H�:���NMυm1�-��)�}��PVc�_�I�=�d�	�u+�d��\3ؼ	&6c���v�@��:�2�բ]��L|l��l��RX�i��9V}����*�6�9���$�x�_|E���eKr/N*�?�T��z�(���m���V+f�w=���T����BӔY���\�E�8y����U����9V��
35m�/�F;��.�Cn���*�ɢ�zǅ҃�Z�r�XlxV65EB    f4bb    2930��r��@�!�@��OY�um����K�����4N��4~���b<6v ��'D���|/�Cv/�H���G�ʮPc���BC�lJWr���q�O����hUWIkx����Ϸ��T�J�Ӛ�nt��<����`��p�r��-ib��qG׋E9��x)��r�wG��Cvjy�۠�k����m��5�����o�@=�f�*i��54�v�����y��ِ��%�4�4^Z��8��
u�G<�z!o(����V�et��u�ڲ@%(�x9"��!@9�(�����UϮ��t�u�e��j]���Ty
�&��@����X�k�xF4O|���Pg��\���v<%���ɊMݤ��ʋ3���vH_t�) M*]�qd�ԇՖ��h���UJ@��bC�'3�����Zz����]��H��p�-5���C�bB�n6�h�+���8����T4i��w��%uX��n���Q����v��Z����(F�G�]��ٜ�l�=�F�V<ɿ�GB	�>����P܇�в�/\�����f�[�S�i�b�=�R�q�nᚳv��Xv"Y
��pon�}o��9k\u���X�f�`#�7}3>4eg%֊�4Hu���,�T�$�>���CW�'��@ %�'�u��ŗ?�(�A!�8t�d�Hs'}�<k�g��~q*-�C�=r䌜��<I簴'I��J�P�7�w�oS��ǆ(�X�S|XI����������.g�^�Z����L�>��*�)eZ�Q�(G�L��j�*H�Y�)�f�J�ĀI�|���� ���}��͟ M�����_]�͉� L��0F'�B������F�zi5	�J�	�EiA��
�턢ڲz�"M�3�E�א��3BS��<����,�c�uOH���t�v%"��-��B5x�*�������t�"�����G�`\Y.�*z���]�ɎL�{"�	�֐T�Z�7�tc?�(�Ow%����e6>S�ID򢻘~��Q)é|�b���Q=U�LCf�G�ڸ\-������|,�ْaԇ��a
����TޫfƄ7�:e��{/d�KH/�nOKx%����	k3eV��(�!/�T?x�ýyuc���G!� �Ns���|%�� ��b8(��A/#�9���j�B���lCܔ���鐖E;�!��Ah�1R&�K��He���&��
H�p�ZEJL��c4��<��-����:�1�B��B3��G�\6����~�&[�a��o\#��`�-f.�ǁ*��d���a6[Ӧ]r�ª�e?J>ʙ[|�}*�ƽ��3�ɦk�qP���@�2�R�I��%2n쌑���&�́�F�^��˚I��5'��ꄅ��R,R�\U�O�;������q���a�B�ҫ� 7��x-���ը�E#ET\߀�u���}vXԈ��%�J��?�R>^��4_�ry2Xv5���A��`�sJ�63�YVD��ȹ�P���6"2�Q�c=��BH�wD$�'h�'��L����@&�`t�G�X#��+��ǢKwH�(c��"�EPЗ��M��'S�Ϸ�2zck���l��� ��/�hA4n�@�ݘ)1z�Ԇ��	�*�X3|?��۫8�j%���N�K�]l��H��'�Q�a#���6�J�i���ѹ��}՘�Ts���q����1��v��?�#�&F-C8.���ڮoO��������M�J�3�8J4�d ��x;����#�#����u��:�5
�B����.�l�h-��hͦ���-�'���\Ê��j�&M��i�Ѯ��ҵt���K`�dJ-٫�J~m�x�~S�S�x�k��wA�鷏 d�&sh~П�8@�f�+��p�L������U���- 	@,�����%�x;@��F��}���<���;b�� kUP�u�Dd���+�,��_P'�����U�ߪ+�H0M�c�m_�8���&
m�����o��m��9���^��N��9��o֦C��p�P�M��7g�� 2�F�v�E��:��4�ؤ'��g����9zT_�#x�#c�_�B��"�l?�I�������1�%UF(��׾,ܵ"�e�ɵ\��S:�
��e��t�t�2��`�Rv:m� "�=O�F���hW
�64�~3��0���\�E�g�#U>������C+~���C*hA���ig��LoiO��� ��lg碰�[C{7V����t������{݌��]%/9ٙ�����/��ѫ���t҈X��^�@ߣ3��J��~��
�K��|~|7hh�������ĔY�qe�%BK5�~�E�RK6�b��A'��u+��ru��Z��͢S�S��4�̾�m,>K�j���c��m�5��{�A,�L�j)��$EX}�:o|JW1P�c����_��3b�r��<)�X}�C�^X�r�g;�2�o����O��x������3���a|Ml���7TggM��9�8�x�o9)�'=:������5�TE��R,򳻔d�`�
.�	>�Ϋ�~G����tQ�mf��)9jDk=�I/$Wi�h4Y�=	���Y\T�6�-U��	�	�9��K��.� E�`��(��ι�"�_.��BP�:d]�5{qF[y���8+��ՁsrK�"x�"w�^W���)��,�-�u��
v$z�XYB1��n��h�J���	,�ZqL�,�Mi��?qGj�.�w�Zg�HT����o5%���~���9��0�hT}�Ug;K�8�h�'���U� ���I��CjSDW�Q���NA��ϑ�yScԋ��ƏŶ!^�{Ѕ1��nꁌz��I�����^/h�|c�	��}�h��m�wu\��*x��N�w1я6�ܧ�P�.� ����1{���#��w����6�Pp���_��տ��,��T�zWi�Dr4d�50�
��
xN�V�oɛ�᫅���^����>�~t3��?��H�`�եqO��M���:�l�H90���07���X�C�q{��rR��o��Y	�E���cQ����#�H�����[e'oH0r��z�(�X�)@5�Ҩl��j$��scy��Q[���f�`�;iK�NUE����Ci��A�+t$�0�:�^� :����]M#�ޚV\���&��a�dA�[A��\[�y�S볧?���ݗ�µ���{O�%/�(^�u>3g����1�Ʈ�q���W�˄���Xƃ�R3�_�J�'e��5D�{�"J���O F��a"r�t�Zi/[�TiQ��v�>T�>�4���$�`D��_�,�Fl	����6��ڈ�"�������Euvmb��B� �X~,�D�J/beQ6!���|ym@�Uf�l�I����ȩ�h���Fzi �'� ��|nw�I�f�~e7��ݒLA�ڏ-� ��pGX��ԟ<>��ֵ2�\^��j�P^�㠓����Y����q�0�e�ݮ�{lp��M�Kj���]mdr��*�CJh����&+��{�'�Q�]bN���0Vt�(�i)�=����sv�0\�n���J=��l�P�f��!��Ja�e鈠鈶Ӂ~�Q��=��Y�Y8��bd�f�,,��dMGa�`O� X �vM�&��hNE�;��A8q���� h��Z��<���A�!�`�ɮqc��&Ԟ���Is�����s|E��W�7?�Twg,�Tc�"�*+��[X���F$_9��q{����>W�6%���/ۋ𑔠�����pXk�2R�i�V$L�s�����Lݝ���X/x�M0y��sSspFz�֏�	�_���lS��`:)]Z�h
�]�;q�^|��l����q�[NZb������(sԕ_ ���#�;�g,D`�p��#!x�ua�"��H{,>`�P��ǚ!��(���Z۱0łMഋI �-��&���run��N��ܜnk0���%�:��-��BA�S%*Swuyj�T��j�Ҵ>�|���+p6�d����J�C�����43��V-���1CI�db��_*+@f��gW++�(w_�M�S�d�p{]���zMI�����N�F��sWu$������s�i�:�=E-��>)�a'��b���L'��%�Rt�*�$o���#������`�w�˺�Y���;�G���B>"�����S` �	���9Ƞ���ls~�~�\��CfX�6^��L%ÿ9 �!��p~U:�,����<O6��PU+��$D���Lţ��Ȅ��w`�.��T��B� Bi-��9Vj��7[@���nX��~"�k;�
���BƳ�'�����1��s��K��ùO�Oy�l	0\զS��I<.ߪ���B,�!ƚt�|r�R+��xy�#O,�n�=��̈́�w
��N2��U4�����y�N�M����	%F$��*���� ���NK�NI���16_���~p�y���hq��Q�ݸ�����`��#L�G����/v5:�	�-��?�VEߌSH��ZxQq�"���7��a��]~`����2PSCzjŘ�?:��ML�������yk��e�8���a�h����m�;�t`TLA=QY��g�fd��q�GU��3�NX#�oJ�֑pQ�.�L��"e�prɑ��=�)�P�"�O|Ev�z��Ct����$��*ܿ��!dz�6�SR��)�<��0�� �*���*J��pBm��i �����BX��`�g4��ƨV��)���b��.Q�fc[|���f�j�Аc�}��&b�%3�"����+Uu���!�Gڍ�-L��NB�.D{��M��,W��	,��%z�|��|���ٱ��f9�\?w��a�AB8 �oN�s�&	)�~m�akVR�/|ڕ�cF�G�̇��R�pt#�M����U�9�P��o��x�x	���(1����NK�a��	��)��}�������l� p	�1>�Hj�l?_�7+h!���y4f�ʤHO������;�~�l+�Z��(.�qQ�l�_��/���QH��OǗ���z�XdtpPb��V�����I�@� ��D�E=r��$i!��'&Z>
u'3 9H�`��?�i�g��Ɖ�.�����Ȫ�x���6�wU2�t�wO� <!JՍ+�KAt\��/Z�WC���*�����4�%�0�1_�C񍹺�����s����:*[">)8F�\�3�`h�~���VT�s�.&9�	H�d��N���,Wñ���s�iH���ܯ?dx?{�)�j��گ[�F�$T^-�����v��F3o���+g�p�cJ��UT��M�1w����ڍ�tQ���
����a���SC7�h�ů�׹{����k?baɗQf��3#d��K��f�#󑳫�o�U�[5�Ռ|P��C�?���m�A!W���6��q� N]���8c5�J,L�/�/�wg� �����֩؟:\;r�R�Ϻ�N��w	��=�:9��V�1z'[�9��$m�nP�Y�0��&h)�`괨��D+�=][c*6�Q��}�(��4S�.���	�����{~�p��Џ.e�K��҆/��_? /aK�p���G���ZQ98;W�w�r�Y�c�F�n:�p��j
�6�ݬ���_Zu��҈�����(N,ْ��h�L �j\���Ν1�6��z����Pb�W����*�I��V6��:d1��s���1g0/?����w�� (�n��Y��B���$��ﳚ�|Y��e��*ԯ�	b�l��fϙ~�]y����$$��]�w`��!U'��}�^;�@X������&��y,8۫9�$� �5��;~���*l�~�U��� ԲD�`�n��.A�#��K =�4��e������s��
�:��z��{��/؀{֚� ��2�k����%+��E���5��n�Lɻ6E6�L$1N�Hf<e��>�H�c�ދt� {�o�h_Z����� .l��HgB�X��A�2|�.-?o���D��an��7���~��ѥ f�8����p���Qe�u�Py7���P!� ��Mj74�h��cYѷ�g�u��h�X6�����d���+/�����(���v�bP���\ʽ>*��Z�=���mV���S1J�&�����s�8us\۫/d�������������!O�ܕJB�׃�+��o���@)��7��L�K�U�ȌB_��^���O�)�|5�ƪW���:�?)M@�C���`l7�FՀ��|)��C�ƤC�T��J�y������TU���c:v�����;gYMC;��e�"�8�H1:�g���(�U�z�ît1͓�����u�)�{������4+U��/.1c˞R��6L���^������ �N\q�a��_�a��6����.��q�r��J1�]rA��'�2���@�.u��N�-���_�ML7�ގ����;�oB叺 �dsԚ���e�iH���90������_i*T/��;@@D66`�Uj7�`��sEZ
_��D{�L{�M����
.o��T�n�	���8��e>Z�\���|M�{R����ٺ��-re��ֻ��-ه��<��L��F1��b�hD�C;�FX 0<>��I�Y9ȓ
g~~H1> A1��N���x�̉up'�NX�J��|�Ȭ1ew��P�z�$n���������
��@��F�
l}Y�� W_��[�\���n��<_pm_}�-Nn�86cӁj�I]OC��e Y���S\H.j\���c��,R��#>��c��x݀̍���M �m·K������c$Y= �l���3������+T�&"I\����@=��dKN�V��_�E�.2,Zka+��\>��1�2325���<R@v_�|��e��p�G2�ؗ�o�DPС. ��u���=��4V�Y˦'v�+ 9�����&�=0_�̫�IkY"v�st�x&vp��%)zE$#�ܹ_z��D����B9�;���8O��%��N�̧���}�������驸+�.��(��O�d�����[d�ى�/�*������.8��%�������m��O��H������>��4@1�YTy}�HF�X,=��v��<|�!_�RF-����W��0Ό�G���S�7��?	����b���p�J�آ'���_w?�/���-�E��]F�mރ_3�몢?Dq�ٙ�/��U:�������|'gG��e�3��c�3���)�+#w�X�{�k�=����i��	�%��uV^����@X��uS�pm*��\�,U�U�C=,�3�c>������v�j��ҡ����9hM|��^3��w�WȩT�Zi�Q4M6s�ķ[T{_�|C�t�eE"�x6�EgK�ϩXg���P�H:6��C��0$�h1�a{������S@��m����q)�<��9�}����j�'[圖<��U�}��T��<y�{,drV�݀[t#;5az���u�����v6��Td��m���8�'-���`� Ѫ����()�v�$2Y��NM��$��M���.s��y
���a�U6��.0��8�T�ZPc��h�S|���ȣ+U;`�q'�!ݫF���XD..��_^�/��4�͟�c=�At���QS9�`&(@21�M��z�F���'aD�G��V,�F>i��_26:K���l�����Z�	.�7��c�Rp��bS�rA�[��F臆�WA�h������"��	�u�_�j[�m���S��*�a.��[���[��A���*u���X��ڹFh��07�T��U�x����K-�X��N�������z�f��ӟ7*UX���V}��/��5cȫY2����׺�dm��������x|5#ao�`� ��+0ZX�����z}[���>���8���L��8��h��*l�M��8���rt����k�{�kQE�l���;��ݷ�n��KK�.L�?��6h�� Acp/.Ҷ��P2غٴ�j��W���E@�Oկ˿!Q�.�fɷ������j3ZI�}FXN����ݛ���T��8	�MQ;I��`{�gt�f&IiK(��g�?M��PEudZ�tBJ��n�w9O9viG�.�d�-
r���EOW����foF��h��)]��K�QntF�"��n��̶/^�z����d
��wX�Y
q&���_��4����ݦ�����V}��� ��q��h��Y~�i�v����WH�|�ָRe�@x�N�X�u��v#����Nd
�I+l��xhE��H)���s��j���^��Βc��2��m���zh��`�DS`%�YS-��r4�j�z-�y`����2]�3*[���E5�WHe��Y�͛Ǧ��O�Ukh.��9~P�5ݓ�̐vM��}5
�?�Ti�/�hmF�r�w�{�,k���E2�)O�)ߨ�O��j�s��ze��X<�ㄙr~���쾵 ]� �BX;�@t��\��P�k&C�u �9�F����B��+}�kܰ�W��	`x�2
c���k�6�[8����Od���4�z��h�[X�q��E�j7���D���~P}i��� �@|��s5j������8B�ZZ�@�}��E����r�DG8X�:2�0�T7�`o����"�%�/��]�����֖�7S���QD^Ў|�͛�4u�>1V��S�l%S^Kh	7'��(�R�����d�Z��ے��d{�Ŏ��'`:%���3,Λ�'P�����:N
�@�k��|���X%=�C",r�����&2�z<Cj!��cR2�Sv�Ez��h��Ӭ�*
��}s8��76u^`$
����f�t��ib�]��b>�Y���4����tM���	���MW��p�_�m8'�H���k�.15�͖��f��<C��|�W���D�z7w����Ry�������2�Mk���e���p�b��*�VW)�J�1 l��r��]�xIAj�a;����W��93c&�! ���k�A�}:����A2�b�T��שr�{��*��"��4�{��p3%CD���
��|��Cg!Y
Y���X�l�撜����w�e>ºw��>��7.}��V���Ĭ<��֐����Ћ)c4n�Sif�F�gð�C+�@�h+�l׋��x	����6�,_�?g���l���
�!vz_HA.+I=V4������#sCt�6!�nU��:�M3����!�8؊h6{(����Ԇs���ҷL��Tx���P��uJ�K M0ў�NE�Ֆg�l�� �z��( D
���ˋ�1N�i�� �����B�BC�h�;z>]�����e����D�%��}�E���x2��^4;(��W�#��ZL�����]n7�R��5�oe�0>�t�8��{>sG#��5�Wݮ�m��'�OH�n�3:j{X4�L,�uu%�T�{����ʚ�=��ǦϽ�{�V���g�ǩߢ6n�^6ql߲��U놺״Y�.U���޴lF�ݱ�I�g�铿c����h�ȭ|�`�ۭ�d�$���4��>Ĺ����ڒ8p��o.}}[h�ޠ��D�ςoj��p�'��?�GQPNԘ��р�Tf�e��s�T5��:�|���.���x�u���F�t�lA���٘Ȃ3j)I�GJ�4�1 ���5��;�P��L�[I��Մ�4��D�-�� �9�8~B��es�Vu:ˉt���&W=RN77��5<{��M`H�+-�� 8~܏���}8�m���Ɲ=j	ε]wv^����x&<�C#� A�5�Ǩ��B�yB
�:�f}�9�{�����0TF +�� �y��\g����b�_uT��׶R>n�gz�0�_N��+��a���j#�}YC����Kqkq�S$�d��%i@�uq��h�Af��"_�&�g��k����~%4���q�&%��67Xн�Å�=�LZ� ��ŉ��\�� ��^>�(��uG��E������]>r���g�F�F�kw��!1�,
�z�+Ե�$SC||Cժ���?㧍M�FN^d�i�@��?��Q���܎��u!��j<��$�������3�����~����,%�\ȼ����/�A���R�\� �rUܶ2�Oї����#b�;�Xy�ƚ��l�j>�����&?�;cnΌ\�8�:-���J�[��\�iᕕ�j5��w]�Nت�nÙ�%���ք���V����)⁭�u֘�V��7y�7~g�W4"����F�i8�Y��U� ��H�>��
]���T�Z9��.�g:0
k��2��W�=M�|37a���Y�Q�q�؈��C4��
���+l�}��J�ڳ}��J�o�����u��ݠ�j�� n�莰m໸l����k���5v��J�ﰡ�T���\������"/;�t`y�
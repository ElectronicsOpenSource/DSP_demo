XlxV65EB    39e8     fc0FS�[���[K#�ߪ q�]��~�zߌ����dBƽ�̄Ff<<��$�T��6��z��e��Jm�;���[%)�W�S|��*u��/��>�����\�u9�q����K�����"��o�d�,nzu�Q��p?m	��
�<�N:�R`Iz#-暽�����|Q��^+��HZKj�������|��V9�J��b��P��q>�K{�ɻhY���7$R�I�쬶��kR�6�\��H�\G����/�a�V��tb9��!�C@h�I$�i���[Mj�<E�Z��7��������+9`�֤%j�ѡJC�bsNr������ W��HSbs��$^�;�z�pn�Lv�\8OVBR(�������e��p�x���3�-�ܵ!�7��o��Z�J�h��#���lI#KD�E���:*�"����n������/0'����ޝ]�3��ڷ9R��=g���-C�.��Y�*����a�'#����X�hz(kW1�CW��E.�;�W���<�!��� ���.��a����ܽ^���H?�i�~���`�9����1lק��k��I_���0�����
3ѲT��9�F����?�>w:�����@U`�Ga�{`
����(4Ce<	𔚣��=6����5���2�J ����
x�Cw�9�J�rF1 0yr�/)O��	��T��F	HV+2a�)�r�X�#52�1�}�A��Km��?��޾u�r��}�8˷��>��^/�H#�0����|��B���Pb��[Δ+�"�^�y�_zUU�¯D՝R��o?�}�"{�m?�£�,̇�� �4H|d!d�RɁ�x-�D�	鹔u�up����!R�X ��l!����$�^�5��<�ԭF���� �e��Ӝ�Y��^�D��{7kd�ak�?�W�D���#~>Y���iD�T�?�������Ym$x��ޔ��>�@������J��T?����g���+)H{\���\���+�r��0���P#m_�!P��^�Xb�>� �Q����5.7 ��Ť�?�ǆ��] ����8F�7'-jn����c�h��]����!N��������l�7����� �s�bt��vw1�{.��n�����_��è�0�����(�1Q����V�Ff�*��Q�����7�@̫Z�_��՜.���=c�?%/b�C<#Y��0�$K��LbR���, ��Z-�?����I�E��l-���ҴSS-h��VL�ۊ�n��0<M���8oh��بsڕ���H��E%�^떵-PGشS�����F"�v�k��$�^UV���#��l���Vr���D[(~���wʈW��AA%e�
{�C��j�ť���@G��a�҈`_W����f�d�_A�݊I��;�X ?ȯJ�:<��)�赣X��()��bԨ�����\Զ��G���k���4_���[��A�,h1:ba�g�'�9.��al�ö�_�ݼ�f���3p4�H޺o~���k�C�J�ƨߜ^��:G����j��C%�T���i��=J��֩Zh��B{�r ��\/P2���}������\�.6���ʠN�������}'��L���ʍ��J�4�(�E�ȭ�UEK�9&RЦ�?0����<(��!`�c�Wߨ���;�b����8���~���E��������9J'թ������Il�g�qϭ��޴�����<�Ֆ���y�N҂�g�!Д�zGW�@@���?d�Ès�(����:{���'-"sc�0J/ذ�UT�,O4\��g�2�q�#.]z�@���H)!j낪�A��q�Zg��W�F��$����e��Jd��I[qˇdQ�!l�W�>W�� �� Iq��i�c�\���藊�H$��#黎�o�\�!�
	���߱���~6ܨ˚أ�]>+��!�8���!�e[~��@�X6��.L����kc+`�f@�'�$.�h&�����1�f��W��aEc|��"� ��`�%V�s*�^�#��W�̗�39��tL02K_�4ń�B�lg_�{Z`��>�����W5�,��\t`g��`�I���g��̣��%�0����E~�(h(YX�hD|�A�B7��G(ͼ�;M$8�zEN��,8fg[-�ﾓH��9w�5�j���&ǳ��َOpEr%�Yfe&�g8қ��co�^x-���I���H	���B�E��Ӆ���0���:)7$��Bm�$�!t9�12��
��5Ӕ`d�+�HSn;�sm�+�a"�����!<����ƛjTa9� S4�&]�ߏ�6��x���������ux<�*�D�f����Eě��nU�o[��z/��˟a�=8�j��l�nw��\#�k��N�&%<��Y��5��w��7Ɏ��F*)��_bk\���XHY=���LB����g�E�����#�u�ź~�(w�L�)7����$u�mAXM��{p&��g���/}u>�9�>�e�$ȏ�jVˈ= ����zJ	o��D�z�
I��mY7��S��g=��iPJ��蜧�q�p�I�v�d�r,���{�X��&��/�X�ۯ7[�����t�؄�\����_��c؀c"�'Z*.�A������и�1�e����r7��g�+�;�N�C��S�'�U��ľ_	�8��$�$N<#F���7���>��.G�8~3��̤,�%�+�b�36�fL�1���^s����d�e@�4�A�hg��b�4�-F�@���Z�:�������1A��U!UL�'`o�o��6~2�ao��@��V��勝�e�~s���d�yV��W�fjư`��Gs�^��n!��_�Y��q<��a�Ǌg�#��x��h �ʫگ�fﯣ���jQ���v!n3?��G@ߏY�t]@dMX��p7X�m8�<�V�B��QEuS/5ρgz��-�4��'���$LǮҁ��,����'��M�(A�c%F���;Ù�Ǜ�1��%8�s����h*>p�Pfk��һOo!{U3�e�`8���M�
��f���\�44�6-�m%�lb�^��6�ɪ������N"��I
���N^���Yp�S8��3����(䨄y^��W �[$�^חw��dxl(��j�Ҋ��g�.��׹�ͻYƮ�7o�Va�-&>��V!inR�{R��\��,ʤ�W�U!�a�=*����C��ۂ�HН��?�G��\w�%ZϣX���G�6a �`�烛�+-�"�U�/M�m���8{�c�M�{ZɄ �G&eî�h�����l��ڵ���Sҁ0�Τ}�s#Vi�P��/� ���1u�OSIh��}<��b�M,z�I"��
��$�����ROV@m&*�Ϧ��n�Xt>2�����T���)&Gn����ߞG��p�u���CN��3�Ya� ۻ��m�@o��6�b�:��z�D�-C�9y��t�k��<�?]E�2�U��@ {�WgkA��sD�#e�p��煉ʭ`t�Ap�T�3��VG����G��@���& �x���1��
I?kM9pt�Ex)�L������MQ�(Ra��Y������n��zZ�V���M������ޑ�j����ި�rS)��L-2Y�yn.��!�Ny42��O?N�����HP�O��wc��ZQ'�ZmΠ�oU"����s��r��됝�,���M�A�ʛ� *��&�!/�c1[�ߛj�tnn?��Q<2V�z��R�8����*�R��<��3�k6-��[�|�Čy��9�1:Zy5x�<��+2���Pj�6���W}��&{kԝ������h��k�D�d�̥�)�Y�bl��L���b�}��� ���E���_�WfKe�<DB���-N�F�f�� 74�+���ׯ;���r�:�g~�4�Bg.T�jT�O���
XlxV65EB    fa00    2eb0�̹-@�vB��F��2������g��v,+Cy2p�8�57|�e�X�tr�AF�X��N�k��T=�d@�U�_����\&Z�n�0�˟>��r�Vβ�Bp�����1��Ÿf$0�����v����g 3~l��_hҥc��+-jl#@�l[�;��չi�x-�T�V,4�Vـ�C2a���)zb����(t
I}�� %�B�g�(`"j��ߠ-:v�?�|�6+�3^^�ZO�RC��N�<�P�ѳ����a;�t��o�xS��T1ۘ �ŕ�߮��?��������Q��E]Γ�r2����5��""��I��t$�R�Q!�e��p�Ș���Z�m��֫��x��k[���[ q��z5��������sǝ*�K����D��݁�7c��2���F�Q쐑�+��"	����U�ZL�o����F@�s��Dߢ�t���w#Q�X�Z����
8�adE\�H���n˸�F}��C˲��PA��`���|��!��S��jx�딿�Ƚ���4����Jj��Ө���v�k�E�#�[���𐅶���?����A�8�]�-�6.]���V|k�([L� �N���`(j��.�/sV¬���y�{�p�hk��ӫ4����؄r�l����it^��^Ż�f�ՀA���`��(ھIj����V�[4���{Mߒ�0ϧ��T�On|' ��U�1���V���s6pO��O�f�K�K�����W��c䉶�6O`k�[�q�cM�Bׅ�7"���ӽL��j��2*�٦4�����֛P��H'�{R����
��dp���DEP���K�_���RU͝�o�~E
l[�S+�jnf�4��B±�1QB�j������mc�7P�3g�d��Pi:8(]�V�ȩj}�E��`�c:��s�jή�^��ЈO��2����}Q�E�r��P�~l�@����`�UjIS���E����U������	�#�b��7Z	v�'ܠA��#��7Z4����#������t �u�i)r5�oBx芮�$(�*:�:�$�t�gu~�C�O�.���0��mP�DD��H�/���	0;G]Z���c�۹�Q�7A�_V�$�k��}�X�����gUC�W���Ļ*�,��#g��`�Y��c��s�s�u�!ϱ⭿����}�1�d�u�S���|7x9�Q��TWC>U�/ӳ��(ͿX�or'��f������.�ې�$���$�������c�"ΐ���W !Ri#���1��t�(�k���\���"�oPu�Eu�)2�jv�hH*���_�I�d/�E?�4W���k�^W�83�+0�Y�^����xȔ��-P�Ee� ��|߃x��1�,�v���o�w�pr)���;VQ7���pv?5}YE�z��[X(��V���34>}��ӈ+�{Q�j�ڏ]���Ҩ��6H�+zK_Hb��J&S�Y^9�@��F<[��.�;���j�S}��Č�*��)�n1�>Xw�%�5��?w��'_� d�+ɰb�*AZf;� �ES�N��U;����~�`%RKj!5��,�(o�1���ɖ�z�f�8w�|T7X�l��v�l�6�E��gx�����i��Z��.[Ȋ��?�d?2�s�?~ۙ���}�U�a�����|T��u����S���]L�;����'���F�^�]�D�
��lE9]9�|bm5��l�S�����%�ww�ѽ�)��I��L�ج%�����ß�\�$ZbЌ9A@ޫ�\��lٜ�d,���Ø���y�?g�D�� M��}쭸��^�%#�"�&2��;`��,��t���qگ7C��]��B�A��"������������}������e*����`�9�t�k4ML��Mu��dH�v%�˪��4��mD���4��~��R�?��]p���e����?A+��׮)B@�{%��	H����E$Uۉ�Q��4����;c���v	����F�S�	z�X�B����G�&���r�Mjg�)r!g���b��tl%�^K���i$!�� ѥ��]�w����(;0w=����	ly=����&��wx'
~^!~���T���&ભ�8i�#���)\K4Vd��ǎ��>���� ߌ���s��vϷ)�Y�(=����W��$���E�C�u��.,��ͷ��ڢ�M�G�yG5y�y�|���qP5���Ui%��pv_��~ �nV(������=�=9� Q4�A:BlP�6	����Wn�"X �W62��aw���}�ipf�J8� �J�svi�r�
;�rG�e��������Hݯ�p�R�"
c�����k\�?�|8�QhM뉵+��<���x���w.-�@���
*/i����6�p2�43��^�.B"�Ƞ�{��U�D��ƫ:�<s'�EG����uAk,�y��U^g'vw�ᵪR�����r�[%��ak+DHl��G�ن+�}%�s.�,5��#�HQ���e��?�aM����\��W�y�_�-(?�A�� �M�CZB�7��L����{��8�%#�t�};[3��!�	�L۹bQm�Q#vդ~%�/i>)�od{�P�~Z����^�j�l�x�8��w��C��!S�yqL���t�~9	F������~+���,d�O������`-���P]�^ЬK3�H��g�n����0*9�o'#i�V�̐�x0�'U��X�ݼBڞ;p܄��������h5ͬinh^�6��$�J1P ���l���"���ν�eգ��V�g;ɲ�<u0��m
1���$@����	����e��ڢ���O� �k������2܊���*��ݷ�W�	�}����+�����Ȅ�Ϊ���f3/�o�L1��AeJ��NF��"��fR	 $ָ�z������l�7���¬�+;���m(��?U~�Ut�Dv�<�D���:5�OMFӻ�_6Mǳ�1��9/ה��d��B�Md��{C����� `�;������K�f#xA�� �K��ֱ�ݻ{��C��T����9㓕Q�,�Dng����/C���P|/��c7:�ry��k�h#4���Vg��a">N��8.�_A-��à!�]���_A��h�1�Nkoڏ��Y����$�Q��|�];N���1�M�N�sz  >j��dl��Ѵ�&bD�:���[���M�Rh���Yg>��A�^�{� ��?`�S�u6������aߣ�&fEB�53]K��Ց_�׋'�ݽ���J�.`<d�*/���ﴽq����f��) 7	׎$l��`\�<��c)�� y���|�9Ɔ'��
�J,{9�H�d,t߉0}���c/K��j-?<ٲ��ucɈ����-s�8��6D8�O/ԡ��b���&���	�0���������
 �:��#=6+o4�ȃ��[U~D}���E���%CA��������%�>�n����E������Jp@ô\=�-!�D�L�Ậ^�a�y��)��O1�b~���-�@�Vc��J@$)6����でi�*�7Iw��Z@�o���~\��.z���O�**,�E/ �C`�<��1U�&���-h��%�ܿ�"A;	Ѫ4��)��#�:@Fj��PK�5r(&l/�M�*��ɟ��0����l�0��ɠNP���* ���qcS��uȿ�?pe�/,9s��{��b��M���e��?ܜĩ@7vJčsA �s[��c�f-������¦�g���L��{�p���:�p!�O����!�ap�Dm7^A�z�ł��Jq)�~bW��4��q���ǻ=�	aTj3���m
��ȏ̀V���ލG]�hjz?�f1|TȆ�N�B���&���3ߋ6����){9o���Lv^8�O�w ]��m����BC�-�Fu���?�X���G��[~�[d"�
i���뚖�O���ӆH����fY �u���+�O>Ƈɉư�q�'=��)Z��F��l�[W�N�*"�:�O�w �Q��p�2��
.TҴ�:����
�կ^��9z�#��9W1��験�}�y�����@�@�,
Ur�G�0���w�"��Tx�~�y����f��E��V��|�$bk������Gi5�&�Zs�aej��K�Jk^H)~:��7N��X~�)�� �;�m؜��g�c�Wʷ�
f�;�әD!��� zI�.�JE��&��t9']�mU��D1KwE�����/5���1�*L}M1�r�t8��f��`���Cl�k�|ZU��?~.�g�D��[g�
���F�奍#�^�j�,c��ځ߲'y7�E���o��evK�`�	4)�t��̸-&:z�ؠ�]�5�f
L��yI�/�ɨ`s��z8W��S��1��&Mx0駼!����\Ä��sN<��c������3��L�h �O|��/��\�j������[@;���⹗���<�w� ��@�'�U��X�����ګݔR@��NL�M�U7���O����O��5�Ǫ���������N���qLW���q��� R�}:C��9��}���ɼx��NYt[$��Д Ζhu��fq=��.?�pAZ#2M��jOZ"��Be�`	`]ʤ�Ts�zfD�E4o��1��$з����H�
0g�3�8[��Λ�v��p�%iJ:U�� E�4�if�.�g�7��Q�b;"�E��̏㈨+I��b��Ñ<7]ku
��KA��:�����E``i��#�::RR�,i��������f��s�Va��V�Y𾹩�\~����0��X�;�"��b�U��:�A\�d��K��eX�p�����tf$�ס�������ۼ�Ș�Ox&��E�Ef�ki"+�%�KƳ<Z#I�Ĩ��6`�'Ɓ��jʞ�&�P��+���;�@�Z��'&X�>?���`|ȘR�E]�팱 �;%��]�9��nu]�bTg�Il���j�0&�f��y|�5� �ĕ&�@��F����Ć�I�9������?9w@����c9W�x��R(5S����R<���O�C�G^X�u���Ze�ʦ�C)���Ò*�+�LZ��F��ٖU��FY��+y�F>~ď�� ���ZsXA�U�j�@f��e�&C�y�g�#6MA0�)�Q�d%�Ve����
u�RKݭ�!޼T�byٷ/wOj)��%�^�p1�b3Lqi���,U�y%�;���7��QCA���-�Kp噱�iI�{˖y�0A�)t��p6�s�ۋ�W��$ڨ}&{v�iB�3bj�+Q[�7p�Sd�����7�45#A)̉l��ؙ|�L��Np]�a�
¦2|^�
<�ۯ�҉��Y��ܺW;t��} �p�� ���=t��3���+n}���єa�J�8�CN���w�_6����F���I�!�*i�0dS�>��7�;�=S�x�:J��
{����ݘ���H������bM�ϝ7��2>�Au�r��FW���gy�k�Z�t#p�-�|��8�!�YX��6�<�b`�?��<���vw&s-����J_�d�PҊ���F+r��h��ʩ�|7n�`��Y �����=�n���{3 ��m4���
���x��)�F�� �K�o @Ò�4��m!
�!+j $�� Y;B�!gB&o�D�WsS:�͛X��,���ٍ�/�x���8hvB�����s?=�S�S���Ne�r�Ֆ�O�E�B�ذ�_yG���Q�������5+�)��Q����ց4��BP��3[2�߯��o�X�N'�m�$1�`Nv�Yh\�rC�ݘ:�a+Ox�+�I9��8��g�Qq�VLkd1�ƀ?)�6"V�.)q�(�����Ϙ�OF���gm�>�6�+}_}�?��y4�T�9ݟЇkR�0=B��~�]F�(��E&��$�w��d
в�w�yul�!T;���{5��� r��~������(`��6�Z�� ��Q�����4���o�Bx�23���/�C��I2�k3Jw��I���E�Ӊ�3)O)?��/�M��Q?�%�i�􎩷���5?����^-.��Y��!��K�8|�3`["6��n�D�z��&�j�4�N�i�����nB���?DՋ* jz$��7�w���Q+��2�[ �m�:3+��Z휸?���������q�%M��X��N��&XG�6N+$�#��4H�T/�%��Z�.E/�>�iF⬿w|�^���Ir���N�v���5���P1�l�cD#��r��	�8H@Ϝ�Z;U�%���`��4�(W4�L��!2��}"l ��OIJմak^`��5�ƯsgF�Z�(!�>J�� s�d+��W�G6�6G�_�
bXs:&Vc/�(I�|0���]���k���.�|=�cF��4��y��t\�Mn����`󧆓y&����M�"�T����+�"g���5jrtY��3���r�j�ӷ��҃����x|ex�z��,��W��C~>���B��Z�H^M�a9�,�8� r���H>�y�q�7�<9�_'�)�:;j2�hl�Z۩]nz�e����L�.��]�;��e���PH��ˑd���g5�6��Wn��]fڢ�O����9��@xa-oY���+�^r/e�0�j�;������ft�$9��dQ}��x|\R�<�[���Z��0e'"%��Tgt �D�om�����`� $=����ZVjo������!�o�X�@�l��?�U�Se��ȃBs�4wL����m���b^�w��4<4�}���Kw�Y�_�W�?<x���Sy�	'â��j�WF�N�1��N�]���PQ��<RlKg���/)&�Y��a��
�钯�۫�y��9pӤ^��\� �q��5��f�_ r�m� H���yB쯒B�ʌP�tc��S�`�H"-��wO^�#�AG��	��f����+��}�4%n�9��8��:����ۂZ���Z��9����@�����B�)�cxk��I�@L�Y��67-4�-(|D
=���9#�C�$��!�e@��T�o [��^\;k�Oc{O�Ǭ�5�|:t��Hu2�H��W2��RH5j0<7����ľ��)�V�1��6���D�W�#��UR��[������%�OG�����:��K�/![����7�����s�K5%y�5���b�����	n:(w$�0u��ᣫxE�f6�	��D���	Z��iE�6
�d�ƣ ����V/�։��wxF�Bg>�凒WƵ��F���I��l\8��U�Y�#�d��^��D�C`P W _#��e�Ѭe�R��og9'c�����;&j�nֺ-L�;����g���N�Yx#Vx5��������,W_
(T�8�n,�Ĉ�L��
6G\Ј��
�:�����	�����Y���`fh?"и.@Ų:W#��<�����4�<te�(M���)cR}�P~2�r�@��`�1^�!01�EE+J�[�H۽p��9A���)A����Ζ��!��A�Z�ހ�f�� �D��r�(�hc�\�D�]� ���j?O{Ƙhۿ���Jtݏh���Pi\��������k.�kW3�7w���ϫs�WB�g�㟅�6����8�"������(֩��HӘa� �p��bD�y�lT,���[��K�$�5��Q����W"�3i�-A�GEߵ���
J���:���zy���xw�S��heY�=����"������"�Na�޸*~]�%,qv��r"~��szs/�q ��'�>k��3G-���%g�%H�9/�9O;X�8Ϛ���KP��@�e�Ex�!�����]��\J�R:|�]$����Ov��<�Y���}����X_�.�Hl��1�O�	rb��1.��*Ͼ���g�����ۑdK�2�3l�����R0coB*~�����c��(���Ū��#�h��}�w�X���w�Դ$�����\>��;�Nh���T�-���2ϖ�?n�-���d�i��{�߲M���/#`�`��ݗ�0֟�E��F�̈́,����C8�n�c��2y{t�
��x�Ĩ�Y�e��G��8�������%.C�ˋ���;:
�.+Ů|*�$E�ʔ3b|D�&*�h��V�oG4	�['<�͛ �":r�qcĞU7*�?�;L�6�8��uOw�%V?�9-.��H僰��3�^{^)�Kc����n�%���*��nb�:�Z1[����LF��2��&�7C�0�ާ��ŠȨ�č�L���/4}�I�5��K���+ih���q`P8�
�#�$^U��R�6#�1��!�#�^^�0�uu���Z�z���Ÿ:H�q%J��ױ�,,�e/v���9n;@���u���#)���v�N��ʛ\\�2���ý����mQ'7�}d�	Y�R{�ׁ�<��s�)r�G�VV��[d��\�󨐕���R�(�'�*RcWFS,��w�#H'� �N��c:4t��	a�c� ��f�	O����}��t^��J-ȇ��=� .Ri�Дb��t6���#�(Ce��)��12|�ړHY���R���sK��i�_4�Q}UfS�����>�٧�U�����~��W*نUa�U8j�4��`7}2��羨k�[°8E��L<�nR�Ȭ��9u�oc��$J0Rl��t�炙%�<1W��FP��Ҝô?jCU(k1�vƑ �P�#1�ZVI�ڰ�3+X��k�cOjlg�����H���3�SD�Fb�'�B}�9jg���t$[�e�Pl��s��Dj�n���>yv��S�?��w-�wfqg��/��,K{�gO:K�a�^�2������sf>rz�E����VB�T�M���Ǉ�=����6�[
=$.�=�Q5x
 �@ɨ���w��y��b���Z���_a{� ���?8gםP�<����d�#T�I���q�~:|#����+mN2ۃ>h{���i:d��^�i����RTUN��WG4�����O�	C���M�(���Kv���:!z��vw���| ��|����y1�2��m��`Wfp�z�=��W9/N���&�x9�P���&3dd���=���z�,K��T���!��<��r=�����׿�5� %Z�k:TND���b��cx���Ii��4�$��0�p���6U'���x��H���2JN��=l�X�N��n�(1�^W�������M�ɡ��Ό��>^�$0Uә�eHoZ����A�ƃ��T@��\����t�zM���jIX:?0�&5��?3�ǻ�g:��ǒ9X��4�wk"�%1h�J��i�!~�;�����M��s�X"+�ض:������?�P�u�p��I��!慞��O��*�ƯB�mTU�tF�R����ȟ�C�7�+�W�Vr}\58+cG�am*���'�,�K���C3ag`A�=���;7CA#����h�E�d3ݽ�f�2w��<T�%lo�|ֈ����t��G�Of��;�I`��}��$TB���$d #
Z���к�گ|i��΁¨�|i��蹀��#�S�SRQ��N�蛍'9vn�pD� ��I[B��/�I����b�~j�gC!�66���I}r�%��(%��:��UP��ޮ���m�:��%�f?pB'��n�ظ��s+��vsxA9�0�O�n�"8tD�[Z�%
������_]����qU�Q���fD�n���>��+�ϴ:q� �ۥ��
f���I���KX(r�j�GA�ԟQr�v	����p6@�y����\�kݼ`S!�	u�n_�Ku�0i��on
��HU&�>�~D^���#����!��<}����;�P}��rE��5�xNNIs率�u�,E�[����o8�T4��A��-0C0��� ���f�`CV{�`@2t���Da�|��2�d�b|���Pr�}�_@�����`舐~�ɭrV{��ؘ�9�WH�(�2,�"�1���mvA��4|( �;�X�q)�u�Q�1΅n���\�<�ѥ�3-G�^�"{��@�޳=6�O��糸j`��Ј�[Uϭl����\���?�FC�"<F
�O]?/b�gL-��Ҋ���!���	�zar�g+uOqј���d`�����놋Vw<i~�9��U��3�8.�D@�x�ތ�01�f��Y�o�_���ƕ=�.�.>�`�;#�//�}�5�q5+����u�k@��ւ��*�Ü���zB���Vf������K��i��;<x�6Mз�yzKaH��6z��8���Z|�0��d�V:ʠmI�#�|^��k�m��	N��ښ�x�+�1��4�;�Z�JS��fh�%�ĸ�L�Gի����^����Ĉڳi	v�0��Fz�*h�������R�A�޽�7�5:O��\Ҝlaq�w�i@�+ϓ+`�c
N3D��}���تH��]�M5t�K��{9GmW��{�^ʓ����A�a8����$�j]��e�xG�͎p�Y�b`u�\��kF����vن�V���j��������o��\�~\������w5���ϒEs>�2�F�F��l'���>�c 骕�a��h���}E�P,���Q�,�7\��?�D+���n �/_d�l}�K�K��P��b^�Y(��Yz��(C������X"֠�tR��i�������j���d����_,I�d�c�c7I� =?��e���{��Il�I����+^�c��^�	Q��M�
��;�M޹�/��K�)��3G6����Iea�f~��ܯ����]g��E�8���!��E��^<)C�U��o0e>�3��ے���x16�����p$�ߖh7�!�ms�#��L� �`<v�D�î<��W:��*av^^�^�������'0�A!�Ϲ�4���u��U��j"�E�L=���gG:߭N���PC���ҩA)|C�1�5]�4]Sl��|�p�+
�B܉}4 ������6�=T���D��e��P��7Bw`�����z��'���W����2M˽�����!gu���)�oWBDf�t3K&b��\5�Is\|�MHE��b�;�)��X�f^߭��9�jv�l��];�
̊S2��,i�R|�w<�z�D�b�^F){2��M�\N�|M�@�����H��2����m^ N�;.��j�%�5($�����'�o2N|ub��	-�慜b��R�"��ȧl�� ��������&[rf��ngJ�h��T�g�z��t|4½�{��<�cA/-�_���ׁ��j����Z4��ܲUj�:�y_,��B������Qn�|�0���}��j=�>�G�Hu��YD�����t���
��9�Mr���|=�(b:��A��V�x'����i<:m�̫�B��t�E���l�����ܮjj�ō�'��Jv�Ѻ(�+��w�5�?�4TM?��/�6W~i�|J:�7@�H�V�7��?䈵��_��+u��a�`�6�XM@S�$��Pi������s"�&�s%h�e���~A������#���w�^֢].��(�6���O����w�%�#$my�b�������=�l�ȧ�#�����*�r�X�Y����tl���
�H�c� 틘y�n�����w�6�t��7;����FY�a�&�' �����$B���
e��.k<^.%�z�g��ɉ��>�2)8�P�E��p?|�*XlxV65EB    fa00    2750��޹F��i�hq?\�8L#++�8 ���56��7,?�|Ž��f���d�F���
Xĕ�%������z�B��s�`�������&�����,� &��}>���X�Obmn�뺿2d�2|Bw�.��6W�! ���흪� � l��2^j7f����1�wS��ߔ�����8x�K��6N%	.(�X����0�m_,*~����?~o�z���eK7�d�Ld��Ӊ`D���`��'�U�7)6���\ƛC���dӃ�|X0��)���T�K�;�G"�}g/�����2�{�P��AJ�������8��p���]����ѐ�<�ؾ�t����8/%J��_��%=`r:N��s� �*���w�K�M�2�� Ni�M�k/;2�>pQ;�֏����	���\������n#D����5]�ʳ�aPˍ�Z�o;F2�{u��������8�9�z����<*p�ia�O���d6��y����.��/�#�7�K�ܝx�@l�v��:D�a钹��&�y� a�h{�k_�\�~��QL&A�-:� ���sd�P�$�<cɓ�j�T�NXIE��!�N��Mxq.!��^���{-=����0�����Cܲ�%�Rw�Ǫ�"OŎ�z#�/�m�q�����dE� � o�Q�ru���ِ��`�,4^�}B��0�A4��k,��S��
���փ���� C<B���ϔ����u?�f��� �lgz��V�SYM�/S��fu�:�W"2��6�����T����CGS�c��W;�p��!�6���i��o�����.s����H�ej�P�I� �1̬��E�H6R��:������$�
䁰�˧|Of�ւ-��oY �'5P��ո�Wq��a��ކ�����^��i�V-}�<�Vb��M�G��jDS#8�<�n�|��}��>mo�:eH�ߢ���2:���lZ�je���H��J��d�W�ǉp���[�I=Z4��م˗�����l.��;V	1�/�G���oL\������O%�0��I�F�.��d��Bj��b�QP�|_!���9�< :��۴R�Ԭ��~�pP��)z29��n�X�W�D��ڈE��Z��6kӏ��m*_��T F��>���J�H��[Z�
��v�� �{�ro?,�.�~@��I�8>�v��*�h/x���*�	$L�5��R��
�*������Y ����U���PX���,n9X�F�{3o;�.)�~&d��/2V�>��@�$1�	�6o	u7+Q�?t;�Jl��;� QH�����Ąi��%�~�>-� �B��cR����Bϧb��ʶ�RW���H Y3Z���/Pe$	���f{9����D!���ݯ6r�I�W�$�t�Z	M� 8�A���!��w�q�1$�6�s�U�S�%���N(H��̖�f8d�����"�	��RQW�Y?7B�F��o���3��xa�񿩄����)l?��VZ�a�PJD����j��Mڍ�}�����u��hĢ<yD'�u�v�"Mu��ɭ?y��$�K
���RH�f8`&�\=��HmG�������XpNؒ= ����������3�ks^C�J;ZN@橜��F�(s��ް�l2z�:�ѡ(���Y��o_4R���R%�5�<����q=L�糮D��Oهjg��������A..�=y�4�t��/\�4 �d��2ɣ`�v���L�H��U	ގ��SV�e��b��yN9�@��+?Ë���$/[XR���(�@jE�����a�@�'��P��wܓҏc����ݏ�2��>��F�@h,�;��%ԋ`���Di�~��wfa�{�"�'�| �tY���wX���/DS57����{����JgU���v#΍����p�A��_=h������ƛܥ���j���D���~������_�}ֈv���aCD 4L�s����f��'5}�mE�l�~h�Cdv���wk%�
���:	����w�����E*T�)�׭�:��ɋ��I���]ݴ�׿��6q��4u��Q��T�tj��TBٚ���>8wH�����S��Z��	�y�ov��Xs�0��C\-Ч�Ѷ*.ϴ���I_#�<3�2
1�«��̣���@9MT�
Q(Ҁ>ͥG#������3_�`׉���Ϻݖ������T#B��J"^�y1��L�>ԋa�>�gA������e����P��2.d4X*?`h�����ڭ��Vɗ�č�3D�KS��=�����G�IQ���k6��Y����\@�b7�;+%7(%P<-����Ԛ�(ަ�@~>�%QWʒ�FpJ�S�L��jTs!��6��<�M�(M��>�"��Ŕ�EaR�1�ix$.Z��0Q!�cw�Ɛ.X�lw.��GLtІh�Ƣ{rCE�a�j%�l��)�ZL��	�<$��Q��̰��Xl��#��4����kd��/�Z����x񨔡�:w�ՐP���;�,M��-K�@�Bӽi�<S��ۃ�T֑Ӕ�m�N#iT�r�/�YO��FѰi̚�����ܡ�lm�iW��Κ�j⏍�Ȇ]\]#0�M��g�k`�8��Bv��0���F�n=��W��'��фpBc�B}������8�#�gF!���w�}�5��?��v+�<�Շ�Mz��}��_A4\o |����������ׅ��,���X_�ʭ��}�z�$���fW%]	 �9�``���������ӵ�Q�/��8����3����^���45O�k�(0�/����e&gB�"�|z��gVL#b����q%ݒ��fH� ���-���eєk���ssi滊ht��0��,��L[�!#��ʣj���l܏�{��x��-W�����1��]�)���vHA�W�ͥX��L��H��K��<��WOt{^�uPվ\#���s���i5Α+�:%[�/�6vQ�Gb��p��i1I�@��-��6����2.շ4T�V?����/Ӱ�������o>�&~Z�`>~��7o��0�(�햓�	�5d���d�p����\��W�l2����&y�Y	\$(� ѳvbVi���cF���\Va�d����6qF�.�+��=��o8��*`�4�R�#W3�dk�Cʞ��<�=��W�f
9�8Үtv�Y�7G�38<���G�4�����&�D8	
�$�V�����}��N� =T��ǫ ���S[�EG�e,G;�Wܽ��C'*M9���̒�0|䀎�ϘC��
�I�'�{2#��O�'Hk���<>�*���u�h�L�q�#����ȁ+����q�Lέ�K[���}1��fSIAu!��X@��F\�T���`�Z�o�(�#C.�i|�}M�ë���5�4� �@^�t����PprF����oϾA���^磒>}q�#�4gL�g�8�m�T�2�âxA�Z���}o�n�XUט��� o��t��Vxt�I%~/�:��FM�JH��1��c�G����l��"jHQ�Cv!��������g?gK�,mW�_/�s����P�/���H�_L��g�wxs �y�Y�+t��MYNA�
)�Ց�J�C�
���@�p�.W��r�[�a��b�Q�����_.Q��hT�$�GY��W�ܡ��*;U��c�X�'��"R<����$C�,���@}�Ic�t�����\a��aÄ�'�en�t�Z"�0`�WU�l�⌮@�$#	$~)��P�m7� �� �fh��1T�b&�L~�U|�6I��!E:�����/؞���M�Ն���q4�(�qP�
�N����$q�"iZ��%�������;`/紨�����%�R��s���G��	Umh�0#E~�rN�΋	ǲ�u�yyw�����'j&��>�v��������!.��n<��|��~f��>�^o�6S��`t��2L��c�&���?�m��։�PQ(֌Ƣ�2�ȝ�ΦL�C*��ݰ���I�-s��uI 5{	n�Fo�j�$������
�O��{eZA��	8���H�F'��ү_+z�g��G�����ތ�#��!m��L��z����!����/�=,v���TN����:ބ 0�� �h� 61�
zPӥ�FfR�[W)���_7O��oa�^���u��:�9޵_T����S�D��a�DOR����K�\�	ѭ���7)� :<a�v��r���a���na"�N�JP�)]�P�E����̏&���\� ���P��	�Er/��c%{�Y����f6_(�k��E} ���jCq����t*�r��s�\Im��/��yv�i�#w�_8Y]���m�����B8�sB�d�}Zjh?�9��C�א���a����-�%�	�YpKEɀ��œW]����% ԸϮ�t( |�ꖗ�?�.��a��p�6;�9�>�����nŭ#���X�� l뵧{��asfYf/
�d��Z"n+�0�
����{��ILh�\���6�k�X8�.�����қh������z/~p�V�y� e��X�p��x�������8���j��M+���jq.F&�?��iL�
3%��+�lg��ѳFdH���v_��y#M��Ьu//���E�TA=l�XJ�qX:�@��}N���T^�$֡��� �hr8Tlz�5��'��:���R���!�_A��}3!�33�ʯT��@��K����Y�j�(,f'����<M�Qk_4Q~۝�T�������?�� (��L��!Ɖ$;�;��=��8P�~�5��V�V�v�x���Jo,�� ��<"ZlAb@$^q�(���I,�sFN��:�n�i�m�B���~(f��S���k bet�>!���t8>��ˈ��~I�|X�������X���Lt7�2�N\�~ᰖ�>'�[+�h���d���X?��fjBg*b������ڴ���OƢ9�?~`�&a��!�\�F�K�#��Ԇ��(f�����A�ف�ܬ�޶�?�w�,��Q2eX�%%�s�����(0��{HT��r;��.1�X0� G��͕f�j���!�R %ｔRS��'_w\� �{��w.š��Cۨ~	=Ȟ::5kcx��ً�+��+�bʞ�Am6�=����al�A�0K(����G5ŶZ��^�-�¾�D(�[t��u�0?F�6�m��!X�R�Ԅh\���*�	M��m��To�)]�+�^Nc�D�:�`���-���Z�k�O{�`�GO�w���xj)��E�a67��P�_�L��M��[n9Ⱥ�-h�4qX%L��	s.7qn �syGx�s���9�esA��OW��Kh�f� �����?�60�#��!u�93�&�횘����O�a�qD>`$��l��E�( ]˅M�Be�?��yϱݥ�X�u�OE:�\]+�
�x��?� ���k ;qr�^>���G+���-���C:�FkT��>4�|l�u��`O֜y��̛	Wg)��
:�:�L�ɠH�lL J>"��|�)*S+�8��Қ8R�+���j��ə-ԟ�	�KKY�O����*�U�#+�"P�o�g�F�������Y�dbB��jgE7��'�S��˨��ϣQK�*O;�l7�x�m���S�B-�~���G*̵�#���X�W� ٽD�_�˜�+����)�6��o���4��j���/J6����5 �]?���E�i}���v��O������,��=����,�E�}u&�R��ǐ���[1j��������!;����1Eo����
��~��D@/�Vq����+���r�j�; ��u�U
�I�~@
��BĶQd$Y�L�#k��:���w��y3��1h����O�$�h/3��
$�Z�)�l63"@-Ӳ�r�c�>�u���8V�mC�e#cK��l��[F�J�z�����.IV� ¯�T9��/�v���-��9�|�m�ct{����*�z�O�c�9v�,8,[�mO���d՟6���P�x�X�#s�q��:�nu�y��\��rH�<j��P�XQ8dK�B�PK\0iD��,�HB͈�}*^x��@� *��8T�����y ġ�S�O����P�������QĈ���������Ǎ�<�ﰬ����?F�k�\Zq*�Ù�X	��Rx�kϩO�����\�?�%]{���ZLQN�!G��"u�[3;8¸IW.�@k�ͧc	�7��dd��]�=0[ ��+͠��;�fi������8�:όK�Q�i����n�Jդ�f:���Q꽖��8�d�6a׏'�[�c��yUP�M�2`c�@m:��"�y�����(fƷa\FҞC��2���g�4���zktwg��!�S�_��t�d"ͿJsaJ�xz����T� ��Ë��V���i���:e��Џ�h-� (�@O�v#c��]4l���w_�=&��ָ�ۏ�o:��z�se5����D2�8�(&���8����첓س�H�Қ���\ُ��+ʄ��>�Y�l�&����.����I)��%������!�E=�2���	�b�4Yk6�G"�E�*����L=CO1#�K��Of�"�F_�C[ ���z��>�l���9��qԠ-�uzY�Dd����4��� 87c¿���*�f��.�^��>�S���P`�X���q�J���(f�Ӏ2�"�s@A�Ж�� ӵ�|huMw����-����9�[��	Y3ktK "O'�
8hP��IK����=-��u�(tlouI������d{9B�8�y�5�D%�,��,8��B �B�"��L�6r_-���	p�=*��^e��֦��-�r�Dd�������02��6h��Qq�Ȑ��b�V�i�&`����h
빧Oݟ��p�V�������ǵ�|�ԯz$�wb>�_� ݡB�;��0�&Ȥ��u ���j�;:*y�@1^�(�.8{�~��?���*]�Q��u{U�S����"�4Re�W�AfZ:k'��W#�#���N�(��%��ĕraNT�L	#��'��5V��}�R܁Ǵ��� ��Q���'�@feF'�C�,/ővS#��<K	�*��m�[Vw2��B`y�Y]TSZ+[�E��GN"zy��{~}��Ͻ7֌����Һ�sZk�=�ֶ�y|W� 
���ͽ�D~���o�IRe�{��K6�o��<ɰ%�Nj�4���}[�z�_������a���q_܈W���FIy�����?���cb!��#��0pm����1�u�� mZ������F �K��}h����<�]߷�RݷWY����(ɗ�x��	@�[	�C����$�9�^����8�������qc�b��f��y:mJ�m�{+ґ'���Qy��i�7�����tj�1�p�ۋ�x��	�W�k<Qx¾��?E${�Wn�f ��&��1%�C���1l�_K����s����Y�t�[\3r�t��^+��He*���C�S
����)@CX�r��\T2ã�*Y��fqɪ�N|O���V3�ek��A�]fL0x��3����mRQ���+;r!�I��\����'�2}U�A���N��x��:sm�s�@;`z���RfNSƵz��.)�9��|�w_���7�0��{s�
�?�O=��2���R�z�cX�uY�<��ԇcՏsΞm-�Ķ��(I<�6y���a~"�h���7�Jh�j��O�uD�h�+8�I�!y�C��K/��-�Û ȕ��=M��"�N��C���r�v��R����U��7��2�uيlO=�]J摶�7�?�)���S_���3�(;���������tu�?������猐��r�\bCf5.~��~�x���s�͉��N�~"�,qc�f��������2�ٝ���ڨz�?�8w!��8<Ŷ~�.��ʅ�i@+��Up��d�z沆����Q�&,�٦,�s��𹻭�հ�cզ%n^K�U��T�&1;I�NF�o��r��n�?�k���0���s��DG��w�y�#=	Z�*��M�!�@T�������Y���A hjSe��������e^�jbZ�,A`1�eaZ��Pp�#G� y5����MeB�.q���������M�Nb�^T��'ۂaXB`ċ�a�Ʊ�g+�I��/3�TFZ��5f�/�&t���C�0�TV�e$�W�w!6��e���/�4/R�J�o�u�lIF�~(��|C�jR�@&U�O� H#Fb�D�տT��2q���J��w~���2�վuȜ�mz�;�z��q�o�(Ex���=���А+��v�*�$�����{Ϟ�'Q9����HM"�0/]+�� <�������8���#�Ʀ/0V\{>�"�^�]��8�J?`px�%Ϻ��,���ě=�]ŧ�\�,�q�ZF�����3�Iq�M�.T�+S���EQ�2uA3
���	�	�]mx����HލY��
T���M�i�,x�?�*z�N+=9M�}t��`*���O.A ���b�D��\��𤡎Ƈ
r����8Mˀ(�H��}Y���X�5����&�����#�bǘ�#i�t�w��H̶|�#��[`�6��k����8=�u�@>�_����(�o�N�h�����x����R�s�=�����60c5�����}��p�й aZ�����-�v�/�ur0Z�*S���-�.�V\7�Dm���Z�\V�fgE��C� ����iy�HE���|�e�/�ʏ�o=�4�v⁀M�����ݸ6�E�1�n�55�+����T�CQ��;��:�Z���Sx�R�`���X�G�W��StExݡ���@0W���*.1��I��R�|��\��XI�f��O�����.+Q���xS�8ի(,�	�l�ŷ��?���|���Ϻ����Όp�_�i�ҚF�KuC/�a ��-���T1E{��&��V.4.8�h�5łh�� ��&����vd�~�E�
K&���и���xG�]tq΀�?�+�������Q���.��b8��qU�M X�Ep�c�gv$xBL\O�p��L[���aw���Sv,>���f��D��,y�#&H�Ec8Sp�ό����tV���0���L��?�Y�&��(�}��Ʊ������'��`-��K-�h
MO[�zl�_ЫL�R:�`�����/��K�Yă��G����\D�ZH˶���n��qG���Gk��A��j)a�l��_�Je�<���u���Pu�eδg\/�Ӣ�����]E�@�v���OB�fZx_.R����9��5�tD]�S�"Z���S s��+H����A��c��B+uK���P�[�����r�x^�/�v�bJrw��c�0�!��=�:K0�{�	�xn2y�[��J�O>cz�i0��u5��G$�����b��;rRk��y=�4^y-q7R_
X�&��pj~�� ��
�6��\��rm���v�p��5��ʣ�54zTvp����;\=�CnL�j���`)`�� y�y��iү J�^�[����}�Z�@V�]s�K��:_ �����P�H����uO�^;��<��o+�Mwt�R��`�nS��j+�J�Dc�C����>�)8q!��9t�]�之��m]�C̨�V����b�r��)�ӌTP����*���5��শ�4z0��:+xV�%c�\��jU�rA�i%j=Z�"��j�S^�D%kv5��\Qk�:-�ɊT��:�`��k�\�Hf����b��U@�	�ϳ��G�$�H�[��������k���n�a@?d<���\�$sr�^)�4!�ź�_3���\�v?Z�Ry��Bf Z�\�6@��!�\}�r̮{�X�b���!y��ہ�/XlxV65EB    3176     ae0�#�
y$�/׹?c�>FM@#�Q�5�ӕǴ�Ivv�t�^�U:0�u���v4"r�X����<ت��n���\Mӛ@��u�-e�5��_�xtȽ!�O���cu�;U��Q��R���F0�����Z�-N�7q�,����T���j��q�BF�%X�,�7������$H,fzI��/X2ן�_��I���@_G��N�k���&l�smׯ�28�8�+�QM���x�
/�C����0��������=�1x�6�}�#��s�.c�� ���V�t�<�xAP ɔ|��:8����j�z����s�\W���O�7c�Խ<��0U(*��!1��ҍ����7u��V��wH�L�}/)�/h��O��-O��{�q5&uKdb����A�OӘ��x�����%��������D(w9.�V�]�qp���A��7P/T9yY���p%�m�5�ж5���;��n��w��h�ֳ�@8鼃E��b�ó�-]hڌ�D����R�	��}��r�c���|9�6bf�h��� ��1�����	-���'����}U؉�߈u�@�B̠����Ά�;=�`ew1��m���+��{@�b��?����	C���x�zY�N��������m��26�.B~X ?(!����y�B����P_'j���a��4�C�pG���wH3PC�">[(]����S�YF1|T��C�? �`J����`���7m�Z�-��)?��0[h{�x.1q��5qr��pTrY��'m�#�&a�p2��%�S5D����Pg�o��V�Ǒ5rgc)t�q�­�a���D�s��
��q@�(m��OFY�g2�j:)i+�܁,�[y�X�&�^��4�6�%��n,��m>��u�d(1b�e
�B!7R�Z)u�̱L4n?v*[pb-"4=��
><���G\kڞ��鈶���G&G��A+0%b��}��n8�EI��6��+���S|��~���[cX�X���Vĭx�P �w���7S�!xм�n+}�?j��s�_�LY��VV�k��ܶ���]�h�����7�|��!�7�~$I��.i+�u�9����k�^���[���bĩ�f4}��Ԗ�b��^=���XJq�t��w���P=������`{��K�	�c�>$%���8����L�_�j�p��W�,�ᔚ
�#�'e��+H"�b�1��Y;��Dˏ�SgL!Ckf�h{@AK�OD���IL��6f�q?
��B�|!@�'�+�|��7A[/D|�/�I���,�~?v��;�����RW�/��c�~C�&��g��dillQ>���E��<��7�C�U3�j���ޭ���`��ιV���ɼ``�(d�'����z<o��d]��W�nȕU`��Y����iK2?�MZ�ع�v|�Z�_���g~��N<�&ڤpmNc^�i2��:&S�ͣ��&з�J��_+@��-G0���`q"Ep��d	m��i"(OP	�iM�]x����]�H"d<\/��ܻ�	% nݭO6�߲�5$��!���@4��p�8��ƥ��1�D�9�L�?��֓����@U�!VD޲��8w�}7��q,�����R� wP>�$�Y(��^8��D���_�<.u��d�E�0���ͦ�N�m2BP�W$��j���B���%lXs�E?���N�{�OT��IV�Ȯ�TxE*��Ƈ?���M�����y#�/���s҅����3�WZ��bH���.�)�H.'Q��[��;P���x�����������5I>���"Q����(�u���smYP<���1�%ٕM᫙�\��X�v��jsɕ��A���=���!�X�m�G���b����:�Ru����C���]�F�hО��#"�Eg`��y���8�$'̀�pQ���������H���}��5f<�.W�9�5fj��g�{rtq|��R�X������ן�A�'���|�.=ܘ�v%�[(	�'",��g�$�����&豕 �a���ijܔ�|O̓*)��D�zH-���^4R�*�]�+��՗Cۇ��I��ȫ
����y�	��!�~BW*N���k��KX��lG�?�	Uֶ4��s�R���P�M f���+�W(^�1,�36��ncF��a*�;��_�rDչ���+8�X6�Zm"��7�D2��֭�D� �,�iy?�yE7�ad��H��9&�Q�|c�ƺ�����Dr�vi���m�}��B�'d�����h�{���W(�'�x�@�ǘ���(�i�f�⚟ �����1�/ Y\��ն�z-p
��q��
����w�^���t��	L�����ɸ��Z%Z�0�
�1l������2T�V? y�<�Oq$��^�CO�H7��f���Z�P�jxCPC�ΌW����!���.|��ף) \��䚦�\�Fv�em�����WNԋ��S�-{�C(�#b�V�y�h���P����7�
����:�U�^{��� h����4��8%��4(����	'%L���N	O�D<�De�ُ��!!���0o�\�����D����������|_���vʳ����D�3Ӹ�)鱤?
�W�{@f��G(�P�����e-fŲr_]|�o5k��<'�4��;qՊ�4&�N+����]��uY�c�T�x�#�~�+U*�o�F2w����Hy��.W�!up�I�3�چ"�{9����Q/Y��7��O��)H�ϧT�#*��F������wx��-d��M
XlxV65EB    1337     790��Tb���ޗ7��-.�!ef�-�W�ߺ8��YUh��D�EY��-��;�zn�ЈȚ(x�Ԛ�ͯQ^>�0ȵ_=�aR����s�c2�*&�m�7z���F��I�-o?P��3˼)����X�2��i�ol�nprw���:-eXWm�$JQfJv�^��q�;��ÛT5����!Il���V[x��zm�o�9�.w��kr<���������Rfim�ޱ�1-�o���eg/^�g�8�����ے��Ow�Y%�=G4��_gd_)7�" �zML��������ݻ���ߗ����u�Q��wqQ��HR��� ���Ф&�F�cI^���s��^����	�@�F�J����"��+��W�����-o���S�v¹_�7�U]ykJ����S�l|�6�%J��Q�v��p�36��/��X���A�j]vpn�EJX��Zf̣����VZ:ɋ���r����vj{�6�=� Ҹ��2�%�CB�Q�����l�T��B��O�/��]��hJ�P��s�������^:Rw��k�̣SȔ����5m�j�:��O��J��%O�{rpA&ع�e�n&�����:\��[�2y��ѝ����(mY�TMa�5'���o�勤S'cW�.��ɻ��J%Ŵ��n[]
P��� �b�*�}	'��a�4�J�Jy���-0�{4���#ȶj�d|����ئ���OG�e�$�_���r˻.eE�1����)ó�׾b���i*��h��?��pK�Be����\DUM�v�z7^kS���k��Q�	��i��g�	ڽ澞��|�t�a���������G'�-��y���4X2���K:���^�ֽ9�i�C ��PP�,��eS~�8�n����ܢ�YЊ��-�X�uNay��F�ZF���!E��3��~T��Ќ�<��۫�h�)���[�n��!�V��ɞ�~wG98n�A����H�G�(}��Y  �c�j� �G���X:��e����/D��{f-���5G���b[Ōp�D���/���Q߽��쫄�����r�z%
���tx� �)���}r�$; �w�-f�/w,&��@�>�V�����`�0�&���p��Dw���W�Ѻ]���ŽUv���L���5�D�K��<�^p��Jh]B������ep|ښ����:���e���U��P˓7V��Ǭ`��U#�&��@�lr�`�fx:�u ��=�V�6�_0��������h�v���v�Uq�����7��g�\����P�|����Q����a��S���8GQ _/;h��k~b�T7H�"�|����Șו1��k�;����|��i5�M�pA�d��ӳ�mj�Kz�,:�5�҇���Po�K2}���S[������:�Bi�j=�#���Ձ}g{;�'���7�6�G�q���o��rq(LaFX_HQ��fv�
�����J��jax �����*��$ˌ�������5�I��3��P ��VU8�6�;˅��aWh�} Sf�Kp����Eowk�UJ�k~f��F�j�������S\\lǌ��i���#ߎM�Ep��J,d��Z� � ����~��-��x
�"�����p���!${i�(
��.��.0%�5�մ\:�_C�Dec���Hi0&��ؑ��Yp8����+���Dq|V����[=Ns�%CR�*!��T�k�S���m�kOs�v���5��HX\ﷱ���G-I��T���U�O��[��k��$
����۠G5�-��9�V���t��>��Wޕ--�������'������W��1\�2���`
��3���#q�, ��1�Z
I�Ug���lǣ��hZ�T�w�\ߊ�AqPj��TF
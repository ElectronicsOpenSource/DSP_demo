XlxV65EB    4036    11b0.�}����p|%�= �5��@��Uy�,;� 2��*�T5Zk�:a�zJv9����,+-��%P��p�TNG!��b�>g�0��@��_� 3S����^�ّ��l*ֻ6k�rG|�K��Gɥ��8GL���� #��ʻ5�Tc)Z%z�j"7:4�?�EY�V$��(�ڶߨ�tϚ�~����_���@tYN��ԩ��ҿEǡ��%��j���^����W	�o��ƿ%�ɦs��
������Q6��Bl��ܧD�a¶Ϊ\=����^;΍YZ��qj��'�i���P��ה���M$������:�CI|��ʤ�9��(啩���ϼJ$��wP[�����`�R���dhxE֢�
$�����-��q����
>FTK�rWh([nN�3
7��c޸Ho��� ��ٸH�ᘼ��Ix`���Ĕ���rv��w�n<�
���]S�u
��!��Ϧ�-��v:��?�A�M���r_�+Z#l[�u�DL�L�A[��-Y%�1����������>A���ȑuoZ8�He�����պ-$�|	z�.1X�G�
}J���@�����e�̓rb��֞	$O,��\JF@��E�p�d�[=Ƴ�bޗN�QL��N�������&�h̓��_�T�v���F�#+�T=o��G�<�b��o���BR�bs[���X����m��%��0ց��إ}��yyq�vn@E��՟ta�OB�Lc~�W-��2��+f����������ìG�
�@��&�i�zhh��3�B����~@�L(dS���#�G.�>��r�0,={��5��.03}܆���'ww~*�ܚ��i5��?�4jmW�m�}��P��|=�O�r6

�A����H-�ͧK�0`ِ�U�*���C<l���Md�ީh�]H��{W0��W�h����,���!��c��~�6|���-=�}�D��laAj�zGi_<7	7���!@������Ӣ��T^dn4]F��e�����e�I7���h���ġ]*m$/a�#�v֐*��������S1�S���&x\^绪H�8�C�,h��Dm���.9+ȹ(����Q�����I.<�==G�xY�ʞ ?�Z)�]b�*��=�W\y���|)MÒ����K�-u��՟���R2 jb'B�|zs���9�uI�PM�E���^�'�s�+r�����N���[
����3v��>��d��a���+��Nj�;������C�8�BjԔ�!�2��V/�^ ���tU.����vၞL��Q��f�B���QiaD��=4ܳ�86q[q#-��*��ũ�&�ɖ��.\�i@:�O�I�i�����c��9sň��D%�ҥ���7E�*k�q�zf�;�	f ��c_R@Z}X��:��O�L���b��?��[��J�����^�	� ���%��Ǔ��͏�2�k2�ƴ
&���y�p��r�Y�:7`��:�ix�(�:Y8��Go����-��}��]����h8Rns�M���V�^���������XlɠmЋБ'4�c�K��AB�׻ �<��������2y��hP��x3�ܮ@��<�<Y~�t�r�4�	��d2a��dX�9s��gp~ح�L��a���,'�ھK�sx��ľTdo��_7f*���oi���&�9��e�c�]�q���X78LF�6�sɓ�y�Y1���4�(�J���-��Z�x�u�%�8�ۿ�H�B�E)�ҫo
d�B�����V<�ͯeR�J/�֭��R��S�&.�zF\Q�x-�y�ʓ�Ȕ�3���F�'����_̆��,Ӕ��p��'�A$��ٌ"��2�ѭS��ş��%����xm|�4��F���
Z�>u�����A��'6h!BK"o��v�&�����u'8��`�����7�qQ�MIД]U�Ɓ9"�}�\�p��w��u���j1�AKl]��*�T\4��9[tR3Bv���&2�շA?N[���R%�\dC��2��jۋl����C����DJ�|3�%'IY)yt�]�$�=�^������b ۂU?��m6֓����l
���K��?���g"(oZ����3�L�����%sG(߾�D ���i=L@)빋v8��0�ߓ �[�>�Q�����E���S-�Yx�l V�Tz;���6�1���^�I>����=�
LY%}��o����]�9�H���_qf��9H��4=�>�3+�n�\m�H,p��ĖR q����]!��
�*>&����)"��tL/���x��;�6�>�z��x����*^K Z��m"s�^Ÿ=��&L�y��}9�X�pj��1LL��#��4�m�����$"�EX��+���FB��7e2S<�@�e���n�;�����l~�>׫)�H�e��c�,O(CV��3C�c{|Mf���C����~Bn_�Gֻ�T(�:���Ѕub�`�j�}���Zc%Љ��TX�4S.��y`���{�5ܮDHRg�(��[���qV��Ej�J�-p������Ԑ7�?�2�$����G������j�/�ݰҧ��BR���?)�"�8��9ib����5Jn��򥣁<������98�2�c��� ?����Z���sk?tQ� �81tŲSǰ��tY�[�E6%H�Z�7�r#�3�$E$Y�
t ��	��7�=��;����g�r9�k�٨��v��'7�rcU`dh� ���6��"Y� LS	��,I��6��P��m�s�]� �����m�M-�	����#�Lﭛ%䘬�7��>��&�0�^�!�ZqZ)�8J�n�)
���2�%�$��4���xH�8���OI��s�x&ҹ,�D ��F`쫎�	G?�R��?@՚@�@�<Z-���S˕1#.���u�;m���7�8֩V���OM {8�@ov�.��%?H}�W�pj�P�di1�	X���U�}�^�/	q���W9M�+uϟf0�7Iax��+���`�6���ａ�.eA��0�gN[�i7���í�?�ct͋��L���Q��D�&�m�OFIH6�N��M�6I�d�@X�u��.`i����[ߑۈ1MS�4.�� ,w�yw�sy��� )b(4/^�ސ>�&1|��T�@�9��_�j �����B0���+OPݧ�J���"�)�T'��O�Y,�B�Y���#�:��d��)beW�+�ȗ�
��6���<��ԭ�F�F9K��cD�U�{����K�z����Z�%]�ռ-Y$�Sj>K).m��U�C����9���N�WLv"8 �-�Uԑpѡ��������4"5�)U�`aȃ�/�b����
]�pr.d��"�o��2~�Ц3LF�-�1P�w��h	�J��P�un�@��^��%��}����QSﯸt�U^�F���]��l�h�vhݡq��d[?��tM�Kq%<��r��U[)�jP�+�[������� B��N��^:׻~�G�]iܾ%:m�>�>@��Ƚ��������:��8���p.���*�7UJ��'w��W��,��z55���nb'b�(���L��u��(��\�Yl^?K�p�_����R�~q�t��1��E�`/>$�J����tFu��8"��l�e�%a��00�?��hݘk.C��n����̵����������ڸ̶�mШ^������ �g��%����i���t�k����o�W�G�L�E7f`�K�劸b�B�}�an�SC��t V��[�\>eF���~��Z/�5/f��<G�AT�r�,@��q��"�s�Jȼ*�*�7�:���eRX��1YcjX���Fjj�sy�`G�1~N|DX)񩁡����!�'l\V'�E�j^mt�L���[��Jh�u����;�p�-���p/L램�,���tސ����7v΂����mѹ{U ��`?��6	��Vq��tP��v����ZWqm����]����r�>���č��"���{_ɱ����̸8j����J���eR�o��%�){+� Y�~�
�H��F�-⳪%~��fo��3���ŸE��iQ��=
p����RFf�r4�T5�^Fc)�O�JƷRg��:��9 ���t��;���<f�t��[������Q�CH�\�dF&.T���W���+��FM��*m�¨����pJ�'���1���;zo��������-�'����$�~���!�]����.������w�>B�3�r�q���(�gYT �έCʼe����b5�������q��.폐R��T��`��KGE��7ȚU�P�����؎%�@�=g�c����\˵��M�4^�7�4,\e;��N� K��@a�uP�TC� ��� /��Aiڢ�y��"� *ǧ��P���pm��3�'cT�e�F�|<�fWa�?�NGm
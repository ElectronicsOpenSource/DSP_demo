XlxV65EB    c680    24f0nRje�]�)�2�GB��U��>�%���ph�6Dv�sq3W��ݮ���ͽ*ͮ�,g�)���BP<[�����{ES�߸�O�S;??�Q���>�j	��.x�5J���I$��?P����J�%Ns��m�	�` f<�I �
QL�A�阱*���7mw���/��]~��*?�%Ĥ��|P�fRi�-XJ�!x���;�Ƨ�`�}���E5�����ȁ��OB�uO���#�b$��X��iS�x,Qm�#�y�`*"v&�kKH�qn������>�v�n&�/m������-�ڱu����L2�;~�Lh?�{I|�f^��|Y�5jC�]��"�bh��lV�6��L��������N|@��e!d�{�m��f�އ��s�'m�&;�&3_���j��_�XQ�R2ݓǋ��k|�Jz ��?S���hH�u��rC�!����0:�
��F�uN^h��~���
�.	��)e��EF�tq�%�2���=T�4��|�@KD��7�Dб���[(�\��j��z��預��͹x��qO"�����77sS�Ĳ�~5)ˣ���.�!oy�ܩ�%� (wT@�B�$/L>dlȺ�;�9�����j��E���7� �� I?M(F��u^���u���
�2��.�ą�B���YG��s�4"�Zg_1�7Ɵ���Jvh�%�<�'f4�'�x�>�)R��cRB	Y�l&r �48�͗L+G��)[=��[��d0�y�<h�O\�	:�2��*.���3���Mˉ�&rϱ�J���{�x�&��-_�g&�]��6�ETSaR�x������BY��R�@���^�B���Dt,"��H�qE�����^b�����W�Ct�;2p;pD�#3��Uqc�J�4����./`��?��p	|����dm�G� �tE%�v���(�*��*�l���	�8���B}C�b���d���@:��?��;�t�	��sqd�B�l��7�|7II��l��A��hE���uU�/�15��H���װ�=:�«���=ϵ��� ��<�{�(����J�)��Ap᜶"d��HI u���jd��+;N.���p��[�;��Q���	p`,�� *��L�@���b������Č�l�jUA��v�l9�FqL�/a�>��[��3��#�fG��&S����ʾ�ز�.��-�bJ���M.�����;�㥶=��݇���/�@���eLk���}S�e�-�mQwDU:���Ľhi}�
-L0�i�dx�9�6�a���	x�]BO����H�8��n�]F�O��0�����I�����΍rY����@�/���L�$GJ�I&�]�Dk�2
A͙�@1z;Y�����1�'��g�3g���5ZO����Pu{�H��(��l;��d��m:������&�D);���z�v�!ێGWL�٣=���e��
	�<�ɒcr��=�e��*��������z��#�<N���H��~nK�wQ	���=��	��Wi�Z��s�d����/��7��?������)֔�r�Y���$:�^1�Ht���8�n�RS�J�ݐ$� �u�&�����G/[�ժ����u>�x[�Eg�v�AÑ����*T�@3o��Dm����p�FF�ɕ��!J�^L��c�Q�F%[9<������&z�0����bk�nU�6k��vPY�V�W9WRmR;���p�G��m$ԏ�j�T�M����^!�8��j�_�������Q:U�M���,���.�;3�¦p�ǏkK� M�ޡ��?�~[��=�Y�8�jlgdpW��rǻ��9A�}�J})�2�){�&��ܿ;���+�&ne*����Q�92�*J&o��R�Q�,L�~�o2Μ�x(�:�%���Y�g�-v��@�@<�e	ب��s'4��(�-ܝv] kz�{L�3k�f"z�{�r�� XB\�������d���}�C��a�{��5b�ɞ	���y+2f0?������|z^�Sى�׃̚��d��\.;��7a_���s�V�Ӊ����"έ�������\ŀi&}LǾk���rⲿ�������5|��X��..H�,	���Q�藢ጡqݛ����1��&��5��q�� [�e����W���M��vk���/����2ڱ쒌���4���&S�������N������h����r��n#V4̑�Ja���P�J�iHQ�Y�J��"D���}�ܑ/a�,�Gs&���ud*�CtY@7��Rsg��NK߯��u9�j��j�\$�{��Dd6E�N9�^A�>�H⦆��i���E�,B���,w��Z���F����7T`�~�֦���j�![��Γ\Y��8Z\� j���)��O>Mv�ϋ1o��G<�8�ų�!��4q	��z�5���c;q �k��ޚ?;���iET`�%�)��,FY]�B�1����������Y��;�0h��~Ef��ө`���8K7
2$��n�������4Bĩ�ä?�ה�p>`K��L)�})�`���{���?��-���N��9�7�<j�ֲ���7}B�1-8ui�=���*�H��"�&���M�
Ɣ��1���1�V�-ګ��}#��l=̜��lI.�31�gn�)u8#ƻ��(��{Ғ:1,\.�tF�K�Xg����C8_D����8��2=
�lG%-w�ܐ�{g��h�,�0�f�,�|/;�^�����Ӌ� m��Y*[��f)B6E"�0
�x�,�h���d�햼%���]&^���V;�`J@:Ɩ�T� ��3��M�?�q H�~YG,p�~۰m}�=Cb�SWν��B��Ӭ�G�����Ɖ[!�p��5�k�4 ('e�,��[�3�k�s��S��J������O�Mڔ��0�m��vN�!�v�޿�mij��V�U)B�"'Nm>F�㶶W�Za��\�hm͐��T������mB�
�Y�?A��W�R:Y���x�ܒ�uA�(�I���.ϙ�Bh�2ʲ������(��&�H�����9K����U�?�1�)4�R�@D�ʘ<w���]��i�vݑAi���|S�r��DEy��,�p��͕=�z2�qxŵ���j�L�f6~�|ĕ�
��+�F�	>�b�iw7X5��=.��FS�G #ő���J��5�r{``Z��ڔX���<��{,H�׽p`�V��L+���A��%}��W8P�@]�-%w�M3&�b0%���B�����?�M�:�W�V�O�|���O vM�����SEE@�DA�7R�q�~�+(&���@�������6�!�(!��������̕�R�T����W1�4A���k�I�/!38���C����<��
ݭS�WE���=��(M����6�
�rBm,�FvZ����	��$/�^di����4Gl��g��]˶
��U�3)�M��[+�9��u;9tZ�i��$c��FC�Q[��n�jQȠ�=Q��K*7����o!F��$�&b��c�{�MR��������AUف᜗~b���|���*��M|���C�gD�������ӈ7e�ѣ�f�	B��6yEB�s��8P�ئO�ݯ����ݶ�����.�8��@���c�����	O�yV���XN'���-�^d��� �}Im����0f&Ә&�k����g�̽�FҨ/޹*k�7�� �ɣ6y�o�Z�C��;���ŠV�i�s S�����"6�V?�_P�DXQP��P&#a�?�lH1���P��^������H�$��)E�/!�*�ȍ�@/�ʕL�zz�Srv`�Gy����x�� ��%���6�a��"n��N�ה��7��^��8��|���W	�1k��3�1tM�r�o���M��\M�j׸��Ó��3���K�1��odm#J(�&���	���\yG\;���;��m��w	�@v��n�g��h�.ˁ�F2ތi�!�	Ծc�&�[�%(��l�(�W@߃x������π]�0J
]#�A�<g�l�2+�L���~����]��"��
� ���j��v�CSa������;�3��`i9	���&~*3�تPK�}��K%�\�1!r����8�Ա�纍I��-���:�Z�祍�g~�f3�x�&D[�vEk��Pۭʠ��6�U��Q�t%�U_�(9��y�F�>�Y]��f�|�O��tO�����@��.+4�LRX��T�y�f�����Z��V#��^����PV�������]�w�aS����~W�:t�t��MX{��.��0X.蜎�����2�P���&����`X ʸ4-.�]h��x���B���Z�=^)ăgC̒)�Da2䲳�]t�8���9*O����v��n��&�j������K��١�U4�F7a��ı���1/��p��>�rJ"?P���!d�g5�:e2I}$ϰQ��ѠN�.CL9@:Ն�k��z5�شj��E��Λ��¡3��]q�p�/����BQ�T��� �4��tq`�ۘ�k���H�L��0���@����g!PѼ���6�S��F��w7F ��5�
�3^=�J�<�{��s4%����D�kkج�����zF�n����ﮭ�%�Kȿa_���֐�j�zKY^��0=J�m<3t͇����MZ�d�
1]����kk~��Wd�8��{�Ss�0M"K��/
�]�G)3t�i⮴@[{G�(����2A��V�4/��h�[���$��oH+�VG�h"��&.�)�*���fVE�ޗ��\R^GBt��k�@w�/B��EbR�f�΄Π��#��ht�>؉);���Յ|�%�ɮ�s����C�Z��������c�ˮ*m3����Ŀ�Ć_�DQ�`���|[�i�,.l}�|���J���V b���4��cCe}g�T��I���,dأ�4�U�&�潞<j���1ĕ_�rZ��GD�.K�M+((��*7χ������}T0�t��K͕C�e�1��,�����!c+'��pg���1M�m��b���^"
kv3�t֐~DD�����Q�BT��S�!��If�JeG}č�g$%_�[��T�7���1)+�X�$������XD�-J��.S��^�L/WU��&�ˁ�9�,��L���0�= ���C�۫0�D����s(ͼ-P�/\My��=+~`_8�h'�y�]�3��L.��Џ\QX<�ѝV�QM���bh�S�H/@�@Y6�'��
M��I ��G�`�Q�j�0���K+�f�vo��ͦ�:=��ɚ(ӯP%�D���
t��Y����OVt������=,&M+r�\;����XV9Y�ӗ��!P�B���}8����xEҕ�K���`����8����':�4��}��tڧ��N��W^C*�,��.N0h�Tj$��E������ ���HB��	 ���>lµ#��%'KU����<N,jr��{�����i�x�܏����hʈ��>j��_![��e.��6k�t�\]���	���x���!�<~�Mb.�~��JMOAI[?�?w`d�w;�f��7NC��kG�}��crrn6#�~��6}ZI�SA����#;z�_�_�Nr�$����%�Vq��52�Jl����7��+{�s3����N��qӬC�-�4�l�Mq���5E�;*��7$S���7�S~��a�-�Q�e�2k��3sW�ځiƽ^�QO�	��9GL�2�ʏ�H�n	���;��l
4I�0}T�=�o� ,$۵�/,��W;bRU�#�����'���z�tv���e�0ʔN�~�ǲ e���*�N�݃�p��3���4�NLb2��(|5�DR.���OTФ1O�Vq�`� s(m��?\d6���5av��M$Gn�&�T����Fy���s,��g�0�8�e��
�8Ml�~�B�wϗ􎄛ڣ#AM��Q����k�]50Fk�H�?����]E"5�}]����o�Y���]xhc��ӡ�a�آ�l��X��>,�< h�=��MF�S�`�Ϛ���u�������h�)o�N�����y�t
`��c���yY���O� ����6/�ꕽ��J�2g�Ի�I�NZ-��fE����izsUտ�����|R&����:�bdW��źl��o���i�*u>sw:�@�$S�`��B>�cq� g�˱�w`n��;l1�z�B�T��j���RBTSW�|�i��R"Q�j�=�����'%ʔ3u����>ϟ.�Iw��blT�bnC����@w:��BW��_����E3�j�p��wm����������c+m�h��Q�ΟR��V���9M%�^�oU��N40Q��%5�ɂb�}mFps��-E���FC��S���#�����6l����|��4fu�$�]L�01vC�����q,�J�"T�~\ 9�?�{����I.#[@����qp��7c�Cy|�:#ۤ���˙��oLi�zNk'�x��Y�p�AwvY��H��������G�d���Ԥ!r��I�u�i���ŬZa� �s�#T�?�J�QV��
���ԅ�l��7]�D��Y!�������E蘁7O��=�QR�zz����z�	y��]#��@ٱ|�X(v�^S�.څ�1��1~!P�CŁЂĉ|��%���w�+�2�UZ��s�q�g���l���;"n,@$v8W��Ra�Q׿�8�3@x9��<e�T귢� {Ժ���*����SmģEњ-]�ߓ#}m����!��*�����g���M��5����OCa±2���� 5��n)O�������7�Fqc�S����cC3\y��v��Q��]���r#����q�,J[����f~MHRa�ίyH�d��O8ѧ�x� Aӎ��N�x�	��K��݂7#|1�DU%ܐ����1HW�)��z߷�y��]
��T�j4.�{z]�Z�Ή76d.���t|��
�'����C�����%U��+X��`�{:�N��h�K�E�#W���N["-F���M��ۈ�̚�9B4F��x}_ t�|�d��̪�&
�y����z�A�k�x�t|�,p7*�\<x �-� �d"����F���5�'g��v!+��1�?ǿ|LFE�l�G��_!��5�ȭ`jz >`ps�8e2w�%���k�1y���B�������K�2��m�gQL^s�{`��G׃�u���sq"�O�ęw�wx�Qj���\�����c��B�֨S����cjb��Y����q+���5�v�֑c����h�5Fc����[��8�ƨ',�\�հj��?�6�D���&u�����h���P��e���!>�-+�Q�EE���8Q���f?7�`#{>��Ѣ95�.�Y�9��2���퇨;�jz�)� !����7n9ȀQ~Đ��(�R��&� �r��#:sw��7o����jPy��X�T���5��s�]��+�*��9�W^mY/i��'�D�h�6��j����r�u��(��-�|f�=���'O̴��/?��N�7���~٥�W��z�ӑ��W@�X�Am��f�ӅhH+�
�<�w#�lw1��>�u���W�8�ڊ���-M�m�����z�w��ᰃFч~������d��WΔ�c��~�mG&�l����Xxl� xi_�'��.l_����4�<7�����~����� �CWOh����Z�)�SĖs���]6�	�W��`)��ڗ�ͯe���`|IYƺ���A �:ܽ�oԙ<�;�Ѱʎ�yq$=c���==���L�e}<`������M>��ty#�1���~�ȦG�����/4w!4��<���6��ư�a.7�u޵Mh��gCl��M&o�A]�ı7��I\.S(x
]?�mW$@��6�+`�O'SU�;S�Q/BG��O���PGl;�d���G5Zk�d�s��q��7��F�w���-� ��s��â2~vR�jx�"?L^(�����v� 4��O
I 4q%z����a�֦jkO�1V]�J����S�z�S8�eǞ��fWmo`m���g��~�|�͌�7$��m���L72�,�2B�4�;�딡�\��?"$fz5�H*B%w�J��$��QJ��+$WPl7
ݫ�#9+�XJ�fĈ���.�em�F�����OYW{3�B�I��R���妚����I)i����L��*��ܔ�;n���
_@̘~�K�k5M���f@�j*��fqz�giFjƛ%US+���������蜉i�c�ZN�I#��W��w�}QFG.��b�	;\}A+��Y�g?����d<1uu����@�H��l�U�Ƈ��.�\'4��V�o# ����1ĭY�:B#���D;b�XD�%�
�n�L[ v��p����H�:�u�������W4!���@��@�y�������C=ѝ)�"���4��:�ܷ��<osa2�7O�|���"�L�\
���ݦ���{LC4���Y�Z0
�ή��\u�i��������4�K�L�;Q�Gw��d�Z��c
����	�:�"L4, W���U;�!���陰�=���4�c����[�k`_3R>p7qj�����}��L�	�_���"���jY�^�9\f]��<�h� �~S%6-I'�H��_����3Ƈ��T��^+��6k0@>8��D�K]I�kqS�o.�y��F�h���1�-�A&���l�T�xO�k��y�fI`��A.�ڹA�򻲈$w�u�8���)��O)�G��C�a
-���b�'�y���K�>?�,��r���+:�i��+�W$�/~�Ō��~d��PfGe�K���I<�y�Ƙu��#��%W���j+:�h3Je_]r��^&(D'�g�S'j�>��f����?���?��T`�)�l�e1*"	<�P^?`���$ٷ���I�v�)�%����`e���u��#��ް=�K�U*rae�MY��$<+�V5l(&�ܠ.�B�pm2��s��]�_�\m��!�~�S��?�?D���2Z�Rn�߮u�W/�\�@g�.]z���[	�IN%����t��u�2��5���$?�II<�PK��É�ׯ��P���/�[Bk�N��y|l��Y��Ju�noҊ}<�f�n��4r��H(~Z���j��Ǫ����,=L�~ q�C��]���@r0>=Lʴ�1%��/�Z/��R��@�8P�d� ��`g��ը]J֟n�ox���^�].1�����,1�"�8�uf;��O���0�
XlxV65EB    1f84     a40������D���b��7IO��+��hr�a�Xֳ�$>6לr+�a:8&^�����S��3��x�P00W����b8,zv����#�d4^ѳ��ڈ㏡@;�kiV��f�g?β�pUʄ[?��`��������W�GQ#�H���U�Q�[�/iXcWh& c�`wx��I)��y�A�&X���&f���^ 	�����6��"<�� ~��N���<ڂB$�|�8?i+�P�/��=�X0P�W���؇�B�S���ߊ���K�!X�{$���S̚ڑz��Yb�
�һ��$�Xv*� �l��3YՄ!��-���Bz!��ѝ)�o� ;��_�H��
��D�(h@4</6n�O H¯�`uhӄq��2eb֚���۴afۚ�Oh�:Θ$8��L+'y����b[,9~��nq��m��b��W[� Fz���k�;��D{j�ֿ[^�h�����l� C~'�k|z}�}:�\ʄY�#�C�ڍ�1�tB/��KU~o�/g�vf�W4(U�>y�'�KSaD�a?��fDP�S�*�I����tZ[�2�5j�a��=���܂�u��`�S���A�v�"7�l�,^�����X��qc�p��9wF�~U�Ue}>����cZ��Y�U�F��k+Di�m��e��8Ń�̝F��λ1�(�Z�c�͙KmB�$�{���5m8�N�؄�>��C�|XXS����1����HD^�԰�ȏx��ߪ)6��s;4��4+f$��y7c�`��<� ͡2�N*,~�M�z��	�����d��0�fr���	]��E�1�֣>���E�s^��'H�0Yϑ~��ᬸ�n�+x1A*2�̀��"t�)F����0 DΥнP�4ԥ_�Qjť�$�k�����۬==�OE�k@AuL�|.��gz�M`���DSˌ���߿w���s����PLl���Z�_N���H�g�J���5���p��`��|��@0-�6z��,I�3,>��K��ʅ�	[�G��* M����\>GxP��hk�p�ذb��Eٓ�&�ܿ�ga�Ǎ�_�����aIy�i贠���s��kp��D����@��2pef�*�]^�w"?t���mi�}ٝ⨙�^���K�}��5?�b�\ �Br9>V�!�W����F_5�}$�����7���Ŭ\DZ�
9z��8�f��%�Y'���@;@�I���E��3��	�Hv�ߋ�K��ݜ�J�r�c�w��&����h�+Xc�����޹���ނ�҂np7^�k�(}#Q��.A�|H.��F[�?�����Gǣ@�"�5���8�G�V6O�m�69��#C��ɐ����m&y=R�_�Γh�[��pN�Q-�e�C�ʻ�M�}L��p�2@oB���R҈C�@dˤ#����G���$ȧ�p�ʒx�C��W��ŋ�Չ�E������\�6�Yʙ�sK� ��6^���F��)@|����F׃�[^D���i_a��gWqn�B�$�Z��U���3?�^����rr�:&4\�[Xr��`4�+�����w�V�����4Q�|?+��%a��^_�T��
�Gk9����{�����&�˸ ��gaWdξ�͛��FK.�a����І�Bd �{h�h�lH슬M���=��P�#l?����cX��������fG}Ъ�Z�E�`�|j�8��d���}Ks��|��f6�$2b��ET��52��(��sI>bo.m1���N�ɿ���#����a��3�E G5��/IU�hK>B��6���l��>	a躨��R��$h����tO�	Еz�1k�Q���i�'��`���p�7���m*κ�<��73�վ?�K�y��q;I�������|�7�q#�j������GĬ��:ґ�8g��*k����6�_$ĞĴ��7��A4?��J���?���$�/J�9p'7ǋf��qC�9/��;�;a�"l3���QS��h(�b�-���Dpo�LXûeQnƸ\[,��32�����9�7����:E�A�VߦH?=$��ҽ�+�'���v,�?�7�ǩ�Z��C%�s��؅�A�a6��q�P| "˟�]�Ur����}5�6f�	�-Sw?+��W��Okh�`�a�ꆓ��,�0e���͞ۦ؜&�85�O���mE��ݹ�����$\�*�5�_��?�F��r{U4�qZ11l�F���5Y9�b�|40���<o�L�a&�m��n�i�����%"��Ku�������5X��9ip�t"m:�P��L���!g23�ƭS���i�d�4�Ra'��y_cq�+4.��OLG5�^A�Q�V�mN�Of���ğ*cU�䀿foss��~��4-6
{���/"����`t��l ,p)K��KPm�G鸃���}��	���y7b�hGV޾@@�^�]ĵ���J���9��LI�C����5��)k`���n��	�`�8�
���%��4a+��D兞pLh�LH�J/�������lz����v� m����RFx0x�[8��
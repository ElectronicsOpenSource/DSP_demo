XlxV65EB    2e55     ce0��E\���lѥ�mN�׾Mo�~��32�C�"���	�|�B �e�$��7�h]F`yytF�'L�[�����'"�W��^O�!�G$���EC" ��0 �ΞҐ�
�R33���51@�S����{\&��b�2�R
���"�+�O�uO�s�_����8汖�+����vaO)��띰
7�^\���#âk���Tr�������S�)m�d|�!z@�Q�e"�f}D����������NkC���D&�sҿ�X����ԩ��y�	Z:Z�ob�F��-���cQ���(|�|��;'ω��,Z��R�2�},N%y��d�a	�����q�N�t��+t��a0����kD �H�ӡ��yqə�E��� ��З�9[�@$���n�S��b5��_.f�n�/�9�n'`�6�?��q'����o����ct�Z���
l�Ә�k����q���q��p�p	�"2v�>�Dq.&���6��)��oe���R��7]�I �"π%v��~4�	��b1������d+O��x�y���te��G	�eb�ܞ�S'�9�O>+얰�;�����j�?����)�%����$`�
Yf*�@/��*D���R�����zH��n��}m�D[��<�$�z�؁"G�ȆS��lU�r�`2aS��uN줬<�2����~y�����!Z/exa�$ӛ�K�=Ǹ�]<-��t16mfaD��mJ�@#L�y��G�i��tJ$cBTc�Xol�S���8�חtʰ[�����0��7���3_E2�Kp����O�#�ש쩲�������z������v���L��/Z�`��f��Mذ^���2C>1Q�Qo�����Y�`"|�F~�����v`MCچ��܊Kʣ'���}�A�)zw�	a��|@�P�/�u�ϵ���w:�$):1�b��%*�������X�wi�D/�X��-H�s�զr�K��Mk�vd<���l���>M	������rWJš��GFd{>2Y�Ө]S,/H�$X�YWNi3����i8&ɍ�Ȧ�6]��%/�`��΂5�S�E�2'g��	99��f�4b��$z!��{B�}��/L0V�/q��P~�&5���B(���X8�PS�I\�ŀAW
������pV�iinva�A�t�W���\���-�u^��X���7r�'%{��S����7rF�-���j�����鸞Rh�^��L��~\I}|9gp��fw�&'(�|u���p0�����S�.3��?%�:�K�۾$�6<Pjߎ� Z�q3��F#}���3�O)�;�ݐ��.f����q�`Є��xSM{j;S"Ya%Ng���{34:�	lugx+}�ɩ�A�
(�{�hK�<���8B��"�8����e���G�;�:�K�K�()_���ZЎ3"��C��۽�0_�ve'�2�|<�E�#�Ĝ�=�W��c{&������o�/<�2��������fS|�I{�>��w���8����f�&�|c���дF[/l�JZA��l�XL9�ǶF��ti5o��9|1��d�K�EV~�#ӋX ��es"3���b�]���rr8<ڼ�� ��^mb����E�♓A����>R�Y�)�{iЙ(yH3�>\�&,06��m%)dd��]*�(RHd&4����
�B���1�ɳ7��-�gI��]k��9Z��Ifd=��P�HFԋ��k��*n��:��I}�(��h�%������VO�M�y��FKG6.E8v8UD���[p�[4�r�24�fH�ǻ�Y�>��Ce��;*"�,�|�AU�D�dd�����:���?��x�w��toz�r�s"���� ���E���z�]����.C	&,^r8{���㸍������N٫3��.�Ϸ����Ҿ�7J(Z!^��^���C!Xe�9����=�P.cY�m�P��AGAZ���r��4�l.8tA�uu,��{���A�Xh��)�ʼv�F�xHEx�P��#tΣ�}h��:d�~ڧ��-c�� �Ə���]�U)�#��~������է�\F����,�����Y��a'ҾU�)��`"��&��m�QĜji�X���d畨��t�5��_~Rr��~�]`v�Hߤ�M��8o(������ �y"	L���f�^ ��ǒ�_(�uj(AêIr]���sī�Hl�' W0�+�< �����G�����dc��;tE� ��{j��^s6���@�����_K���y���A��<7�E��h�8
�N���ۤ17�|���E-z?��%��_�P�� rb�g�7%2�S�;��$fEX��O-[r��sW��糫�q3Ff��b�ipˈ�5{���Ԧw��u	 I��3������)ѧ0�A�պnP��1w9��p��E3'�J��l�� �����dF����͛����x��;�5��f�_!�6k�h T����"�����]��4#�����Je|���vޫ G�6q釓�}Ň�E���;���\�W�z�=���,�#��!}@��9�p��_�ґ��ub`+�f�	BI@���l\v�q�t�0���S�?	Bmڑ�?�t�M� �a4�Ӆ�x��ᄇ*<98j�֣������5'7k" �vy�&ֿ��p����I�'m>cź<=(��_�W�1���i=�-�jA@ơ�|*�=�e#��>�(#{��ڧ�iw��_`4v��m���M���G[~�'�|��c8b�/���S��;�gq�a&V�b�RJ �$� ���!ɰ��_����itc?Q�(�r���1d�I!�Y����L"ȎD���D��Cn_��X����НX��N�Z�	w�˜q"���D�j�P,j��Ej6���)`��@�]�璨�Rc��(o�.*p�?��y�������ȏ�%���@nX����ꢀ.��+Z���m �m�q�A)d\<]K���L�5Tõ��d��$��Z�.�s���]��g��<����v�Q^����00�b�΀,���;㝤�� ����S�)�V�]T<u�Y���C�X��kA["Q>Xkv.���D�6д/;��K4#��ˋ�]_~�@����u�>��hu�\*I`��H���f��N����e���uv�r��@�~K�ANaA;='#M�PU�S7e��XN��eu^@Ȯ�Hy(��d�xI�Y��6Bc��U���ش[=���L�I$��o'��Q1F�
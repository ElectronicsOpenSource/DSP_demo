XlxV65EB    2b7a     b70Q�Q�	�Q$#h�R\���&��{x*��y����r�L��.ٖ�:�$��y�j� �~��]���C�cz(�2�e9�m�a^^��ҧ.B-��,FO;�utd{FdĚ��Ukw�e��iP�P��۾ӌ���p�C��2��ͻ�czƛ2f�ҋ��"��z:�+�^M'�<���D��`�6�#��Q5�h��$��3>��F�b�}#��;��G��I�e��0���.����3i�p������\�y�y�[�_g�	^���2ξ��!��pT��1"��8��N���F�����FB����=��yC4vՋ�~��֦S��I����QN}��z���m	Gl��=p(�)Uc��)�(?`���zJ\��C.���� چ�/�09��M$�����<Z����F=�.�:�z�X���w�=03L���o��*�y��������1i��h���u���Q8��Lu95�!�N��L��h����և���q�q�����]��)���Ҿge�a)Rg�Pyn��������)�E�]u>��Jj�e�(�X/�#l���Xg�g��E�������O��Z�u����z}i���h1"�����g��B��x�	�+9�z�޺�y[�����({9  g�%1\�61�F��o��W8u����Q"�Yi.׼i��<Z��̎oeH�y��e�.H;1��kRX�Rm~#�C�5�i��8}`�>Z���t�ج��W�����S�+�ˢmZ�B`��J5e&����ɓcÔS���􄽳m0��oV��b��L�E�֤��t���/o)�B/Ɣe@@?��}��^�$���(�$љ��e�P��|8�픕�z�1;��<�졁��t���"�����M�1��ݩN[�|�Ξ��
U�E�"�x�R׿�c�m���4] �ʧ>4��rJף���l�FJK��O5��1�[�xt�8�Q��n�vq�Q[��ۚr�\N�޻ޥ�7n�v�/��k+W%���\��u�޳ؿ���C �#{cK
"�!!fg}7�(�TQ������ʆ�?5�P7/�����{RL���Q	x`�5ō�v�F���>'�fV=�mBl�W}�H��_?������!�y|_Y�K}�ˀx_�ȺŅ����z�?���.�����zGp"g1+��L�j��S��ո�<t�P
�7�!6��8ܤ��S�3��T����mj@����b��?P�.�ꗏ�­�!�J�&NW"p���+ԓxX����|35-b��=�o������"�%�c=���'�wI���r9u��M x��y���Ӎ�����ɫ�&�m7Qj�0��C�!����!��`���?�L;�>(.��F4�+�to�L�1��蹨W�� �a�1�!S�U�ݔ���ً.z~)oZ�K��� f.�)N�?]Ϡv��_mL�h�s�N�m+�S=I��"gs3���Q(�f-�zv��O��v�z*�꟏$����aR��L��-7"���y�i��׵����/R�@먕��-�y����e2�K]1���y��k��&&���zY��r7�G�T�79����(5�v"&����,Y�_iFQ� !��$�ĚV�n,��m�f�z²][}�ݿ��o�)�ɣQ~K�ynoCfK	��2���;����	c��E��%L�����H�뚗�
���`�n�ll�@i�uTB���A��t���}l���br����i�[\��S��S!,X�O-�|D�{0JN3�����7��(��2�jz~���A���rN9`���z;��auxՂ����B��I�3�3��Q�m�t�Y������}�O�����L;��f�8Dͩ�1�,o��}h-1�t������ڛA�w���]dǕ}](�״�p�M��)2Y:�I�$r�V�P-(��R0���$�� ��|�o5����=�����i��H��EB�����"!i�������
�dw�м��"i�a��8�t˔��{a�{<�3j�U���hw�-n6�]&p��M��=ث�1�I�i�\k@�io�of50�+�:�i��1�ȹ���C$��V��.�6[T&�3M;m��\1֦���m����3�$�U9��eف��8���u2��!����%M��p2-��z����(%�)�.T��lѬP���3����Ӯ�L;��d��4�1�>u��	��*�ڌÒXƱ3�e~�]*-b�I���V~G'߶
l��ڪ�#{hT?�M�鵟��$S�_����ן��3prL���Ŕ�4��wFى����i;�ՙ�#0r�ܔ�5���{W1n�D��`�r*1�fJ	����<��2>�~W�j����=�w��M1���,����TF#�u�*�tY��a,�Z��j���1\CD�6���$�eU��a�R��㫥�i7�`R��Q:-�;6��T�4�c��G�LTv�ݲ����d(�s 8{�_�-y�E�r�r�t�
���������Sۘ4��>���z��3�G
[��|�ذ򐨔���P�'�G8�/��C�Bi�	D�/�e�h΃aa�i�׽��g-}�+�/�a�a�u8V(�� �?=_T�pS}��B��HiD��ܟl�>FC�k�	��9���H�ԟ�Bw3��g�7/����38�+���u�}�0
G���SSu��s��!�n]p�_��g��%^���V�NFq��r�h�������@x��O�*���=֌��	(��ݫ�-#172/�צ�v�r�,=���,�h�§q�^> ��Q����-��Ѡ��zA��A`��[j�(N!%�=J�Ark�)ư�-�?M���J����_\X�45��q,M\0tg�ǥJ
�F�k*T����Wg��-I'���e7�YN
XlxV65EB    fa00    2d80y
�X6�r#�7�k��Ǎ��P�2Wޔ!�[��|W͉��&m���7�Q��tr猸8���`��K���ewX�jS�C 3�Z�0���<���QM������ ��MN����ݛ�cZ����O�)d����g-'�I���m�=dmqo����&}���Ϳ���!@��('!(Ma�]�0�ّE�`����Ap�/"N�,\-�K�7G�X+�d�s�Gn�f�;�_�Bg&q
Z���ϗb��ä���fy螏5����Q�]��`�t����OI�w�j��1��u�X}��+fgdT��zB-�.�ha��1�g-Mpmv�A����((F�U�K����/�r��u`A
A��%4��k����Qx�(�Q1��b-��w�WO��-�{���P*#$,;�,��ԅ�"������a
��{ ���7�$�<�S��$�	���Ϸ�{���Q�����S�aϥ��C�
bN#�8hԝ���~����3
#�]x����X����M�e����ㆠ�|�Z�l�O.3�9�a���IT;\���<�0Q0��]t�/L!���nU+.��CA�y8|8�B=���Y��^��U�Vs�'��e԰�p)��,�7&���)Rf�����\��1G�244:�ʭ��j�q�0���\^<�*�
���z�Ow!f����d�����C�?�����Y��`�� ՗W�#���l] bz��Io��(鮜ҿ�t�/"﷡kz����l㚋,3��L}a¿	�2.��O��;�#���)�7��^ �~�D�Eaz��j�z}(�騁g���/gJ*��Ӫ�{r�� 䰙�"�R\��Gi�lY�t���? �b$
���P��l�۴q<�77y5eu�2Č:ʬ��DѶS�:ҹ�e"86Qҡ~{OB���+�4i�V��-�Uu�9D�	b�c����2^m%����(����;��冬�rS�J��}�������<f���p$h�ȁ��$��|�Һݏ)�dBL!���dg�@��IO��OP��(SrS�/��n�/p9�#G�}��������xz�2�����썧�)���KO�Y�E]]q�y�̬�W���LޖrdR�X���l�M� p�?�K_�{���zJ���w���I��(P��Hq��d�����pq�%
9ԇ���$���<���(Y�#��RR�'3\!�"yiF�O��:p�P�n3��t�RM	eS��%W��'�ɧ��Z��*�ωbm����|u���&V8cfF���Sœ,շ�,pI$^��@Z+���������py��H�!�3iJ9�kdq����f���Wﾅ�<�㮜�)?���Sw�l��t�Ks��}���e�ӊ���n�����I���LW�o�d���ǣ�x�����į!CH�G��ڰjH��W�e�zp��(���n�0��NA�\��6��k��g�I��|&�,{�B���y���߇7���I�O�R�PVc��Z�?��_�P���'���8u��U��w�upv����ɨ�_A��6pV^��^J��"�P7����k�*xt��!�� _\e\q�����j�\�ۭg��+=�6�M��e������|C�mٝ�����8٭�r�O-���U-��~��Lϱ>�^	�W�����{ͤPD�s�q2 ��S���%�rY_�/	��T!�u�'���yvh�������#@�N	��������.�]�ܳfr`��8��n�^�c��b��k�a��6���W�����M5�F�J���@��j���̴/�kpV�B��!�y�0V��uSw,�
-��C�cTߑDa�ȯQ��z%� ��{�C��3���������&zg�[���(B�M��;/�l�l�]-���#V���OP����[%ST0�e�/� h���
w��^Iz�= G?^U|�/��q����Q\�1Q���8�dz,�����k���_���5�w�YY52,�
�9I�G�*,gIG��T毶^V���xh�q�Ptw�F�l+dw��� LB�w��S`Y?�e��B�~7�C����kq�}sŞF�qye
-���ϦOb.�g��¨BR̋w%�1~E���d��;RG($�j2�_K���z�gޏ'����4�XÛ��}�Sw���vdd� ���M�q�#^Oҡ�A(��9L��Ȑy$7ז?��Y�r�����*9�S{샃��j�g{;���'>�j�B�D������"�ϛ2J�GLV�C4���Z�}�ww�z��Z�~�E�Y�޿"��>��Y�N�0u��0�4�Cj��|~��g�W(7�w���G*7/��<���6����Db��aN��^m�s�8ӣj�ll��H1.�-W���߹8*���*J�(��+�'H-{|��l�*���? ��o�H������\��^�M8Kx������>����4W�T�������G0�(;|MM�O��<e!��h�s�]�~�7�3��5d>������)d���h9$�`����gE�,#��0��'l�t=���qѿ�k���/�"��� 	:���$��M����4������[�"��'B��Χ4ς6W�̈��t�e�sH��(
���j�_�pUN�\��Þ"(��&��d�cDo��|OCR�U�	%Zx(�~(|��}-ʶ~Q���׈̉�QWE���Z�
�mf^��Џ9���xC�\�Ïd�������Ə#�X4����ȲO:+uk<д|/�������	�{��!Iwޓ%�PF\���� )�`��||��I��(��f��rٸ[Y)�V3�<��"e�
� �3���M�&��f�uX�T��`%|���p��t�l-��:%Π���6fȒ�x�Mw���]P� v>�e��xnC�I����'��s�9�ӕ�>����nOԂ	�f�&�6��BI�f�`A�T908�w�o ~�M�|��F��_�x�j���Z���m�g�G���}኉P�p�"�i�)��'h�O-��9���������9�	64D}��8��~��,GTD����Ĵt`��	�1N�RN.��D6[>��]G�*Uf^����Uj(�+��P�����<�6j*�����EL�Y\��<���YvT�A�!�نa,����8���Kϕ�	�T����k̘V�)Z�s���VU�(�f���y�,�^�:����)ƿ�z��A�(���xp�������;glE��MG�C�����Kelj�*��z&����#���ۈ�-0�>JT{�$sՑ#DF������.>=�t�O�Ww?��#Q`����d\�[�É��}�Z}�Vi���
���b��:���m��;��"뼀�;g-#���#
2v��4�!��;N[2,-�m� /د��z��_'m��{uP� �������T&�=�T�˜8���ǽi��%�������r��~����\d?xգ��$�p� �q�"(M�dZ��Xٿ�����*l;����]CC����������ˬ� �ݚ<�7�>&Y~r$����>0�hM��٬�x��g�%�I�	ݢ�$�1n�S�W�y�e<�"��Ń�>*d����AB����5ʀ�;@�v�1[�rO m|�����e7�L͔KZ�x=��}���}�p�F���}���2R����˱�t���� ��*�:��\�, 8ӹ}� ����CoDԄY%K�A,NGC%*�'	�t#��Q�r�d���lx���K��@شl7]]\�����g»�Z��r��2lH���1��Ԓ'ڐ�4���kj��<&��}|$����j�A�s���%tDS}���%H��f�dX�8+����lW�bX� �'H�z�k���l]�t�pY1��`.D�ӹ��;�[z$�(|*̩1u��@0�B�fӶ�w��pc,YX�Z8M�H,�L�k���9Sv|����2a� ���H�;�
���H1RTv��t�В�}�#�|����;� �;@API�y��� �޴ܤ,�}>#.e4��Ǯ���R`~�_ď$��8ǩ
��xIbÄ:�B��*s�;c���-���1��p�)b�Q��+���xT�RE{☑E倚��aO���i�G�����G���d��U+D{��$�� ������W��Yk'�r��W1+/ض���:\�O���an+�^g�*���~N液����=eu8\�j)�lR F1<���'��-j����~����=e�@��j?�hˁK���#`��J��� ���S����� �3|�+_75�2��}܅�j��r�T^fb�W���e��4����NT�6̨��I{�å�`N� �s�D�S7��<`0;얎�ИH%��%��~|�%C���ө��p�� �^K߷��r�a�JJ:V?��_e7��2�n��`�QLZ��/M:i\|�Nn��@��u�;�L����3D����	����-#{�s�"��^�r�
g�}���UV taF�_ǫ`�,�A��%��aQ����e���!�1A��s���������s�W~�S�?�^z|�\wAۀߐ��ܣ�[�FvβJ�9�U���+a�Iz@����dg�]�߱�08��Ĉ+F� ߄7�@Vh�?K�Y��1�*�rZ!)m�g;��wNޖq��v��+��#�)&� ��?Qf�僕 {yr:%B!,�f�K*�0��E�d��*y���s��6����t�U��w���$��`{����>X���h/=gC��T_�qT�j�\l)i��S��X�uPai��O���mn��T�uo�/�j�Y	$���.���d[#��`��p
��]�g*��>+/��Yf\�&pZVIT�<��"ڑjz���\�o߉�m�Ɉ��$	\oN���&�Y^�B�@�_�@G�h�Ԃ/}qH�TǛ:���h��RZ^��9��$/)@�8B���+Ǡ������n��!Ah6�Pb>OG�60��\*@̔���r���LK��m}�q��`��sz��#{��a��R�c�r뻓���;�b��
h-��࠯���6�wS����h�G�82�w�B�'Fc��4���[�%�a���\���u��O$ Bl3�#Y�I4w�t�O�!I���w�u|L O��3jV���e�N��f�B�YU} ���f�w	��X�)�7�rh1m6'M�p�@���/�y�L�;v�!)�I�b�.8�(��0{ryDXs�l$u�S9�m�Ev��E��m��+Cy���ӕ�����g�+	���[�a%c����鵶�'^�8å!>]'�aM`T���6�������,�Gm
���Ҹ�,ĸ�b,�)���t�uP豞(yI��o
�-�h�)�0~n��M�į�#�ڑ�o�5�y�a���V	���B��c��/6�ȑ���m��t i�|��:o| -kA���ֶv���9��8X1P�T�u�:1q�=S�r�l�@�&�]`�Q�.��^���j 9��W���e{��?��0-���-�U��].x�,���"��ǯ<����;r�����v��
��N�c)77�M����b�UW��H�&�3�}>��ha�;s����x�1W�5hV�@G?��ĎG1x}xY� ;
��%k�%o�(Z�f?��	�~�j�T�Q��~���Y��'���N�h&X�� �q�ZM�,��	~&k<�a6u��N"�+�6�"e�d$!HB�~��LHw�zP-��v�
E���}�2lUN��^Y���8��AF�G�A�Iݝ �2�K1 �@����Rpg^�c�ωLw@��s��x�h�_4ߧ�\>�^������l?M�*;�8m?�q�:�Ї���������;�/��'���';����k��xz�h_eÕ?(=
{ZVʰa��4���i� ��l���@�*�3i˪���7'��W�� ���GB:��F��F��D��~l7=}l�{sU�C��(�՟偟w���Ǻ��ᆉ�Ɗ}�6�_�^���`2�3�1D��4�U���'�����8
��"�DBQv�\��.qJ'�::(v[���>7�iDw�h�4g����&*�Q�Fhf9.������1�0x(�����}=]��G�=�ok�:�ۗ]8v�Ht�BJ`���',�hӳX'�iT#><�\���-Q<3U�a�C�=$(�'��7d�����3�6Zց
���2f1)Щ8�K�()�!4�|�����c�_$9�`)�HU2��l@�f)0ącSdX,@���m�,:�XpF���:���ٜ�쌗�`��2͌���p�;�I6� �'�}.����=0
`�0�k��t"�à���l�ŉ�[fO�k7+sD�~J�pȒr<?z@eB�&���,���4�[v���X�r�6��)s��[E��,��ݨ{L�&�ȡ]r�A��U�Y�� Y���hRN�a���X��hd��ŐӶ娮���hcB��j��f?�-c���=�����.y���
��|��)����v*�i4����c�O�8������%����4 ����-�H]2���.�������I����K�F��D"3�:�[�F^�3i"6u��v��(c{8���P ��@8k�55������AU�V%�b{P��}+a�&�]Yd x����-��Ե���	)t��>7�.�xm���N9��W�(� ]X�׀�a󨏜���� P�9Pe���Y�7���"�M�&��2��p��U���=��w�B� �Q�-�{�<����V��j��QvS�#�D��}�6�$�K
S5:~~d���g<���p�R�}�7#���㗾i��9���ýB��ΆK�n*��ߤJ8��\��b����6�&��+���w�%��{�J�v�Y���&���PR��K{o� �%J`�^�Hݹ���&.78UZ�>wu:6=aݽn�{�\��"y[^�N��b7�r(���TK2P��:�?Y)�P2m� �b`����p��}�JG���1��O�ջ��TmS�}�rx�M�2��wM/C4�o�Cg8��TYݤ�@��*kL�/�Z^�M��b��\E�0��׍ˎ�g��|��.��}>�xhn�75i�H���m�A:p�1:�%��/)�����#��4��*GT@QV��O��=4�]��-�e ��� �y_	aW�>$ݫqP핬5Q��<QSѲ ?ʇ�L�ȡ�K���T�Q��F��gzX��7š��	�(уi0�yW����P�^R$�d�Z$�q�T�Z)sM��J���=캵[fc�2�r2�讆$@d�	��+zk��o���5��+�8$��f]ΰ �E5H�Ծ]�]��E
�rk���������{ޫ��觻Y迆%��GYL��t����B"L2q��v�\���Y-�)�.�X����3&�QϪ	�u*l��b�K-�-����%K��N@T�@������c�&x^v�{��w���}ltX��\y �PZi����y������ɑD��"~��#ŉw������Ku7K��A9�70�p�mD�#E���Ҷ,C��DL5�0}O���uͶ��5$b�8�S���m6�@��[�m�-m��L6Z�ye�/ꋌ�T��JǙO=�m �t�x��ߟIK8\��~�v7����+obXy��冲������!��eP��-�1H��.B[��)v�q)4\�3��Emm2�� �S��P�f=�ut��!��}�YMP�"���2�G/.�й���L��t���ҋӀ$��Zy��_\�{(��S	2�����v����d��x5��ι�z���kJ��b��-�Z�&4�ԥ\b�aCx}9�G���6���I|�u�t�8�1��7Or�����)X宮���m]X�\{^�Rǎ@��s �B��<Z��)v��s���S��X�d�j��ۄ�m�}�)"�]ߝ�d�Fp��I݇<�l��?�u��=�/j��&R��xx��q]d�g�TFX��ClCp�q�'g��.�0V����N{�;��(�PI��~~� ��w��M:�LR橔y���0H���#��WJ�a����:�Ust�c�c�}��d1��o��	^~��!��as�*��{�{�a]3����Ė���#{���켆�h�<R�tG I���G����g����̠*rmN��x
D��ƊiH޵fޮ�E��0�;��._g�Q�,"�h_|^pC�$gBuy>�e�e���Х)�,T������sp�n�!�\��e��B�a�{��1T����Gף�$��\����ޗ�n��e�'�K�XW�6F	G��n��c���R�y��P'=%"�\j!�[�	�N^�K{��I8�,aRo���\7�k�>x�s��Qͩ�ƃ��C03z��b�	�?��j!�8gB�9�;:�A��8F��Q���� �3��h�/+x�'}X	?��=C"�&SS�ߔ5qfJ���߹�3ɑF&��zD�����x:{���>>�O���_a �.���1�����bÜ��!	�����]�dk����h1u���{��Z7>u"	 ���H�U�ΆS��;�<���#��ESF;A����W0��Th��3�<�@���3��+���֨5	"�u�Z��������������bi��pfM葵T��uy¤��͞�6s���	yw7Ӏ�G�1;Z^s���������ɠ�ht�`�ӣ�J���-������EL!��1�^$����1�	�r����X�o&��Y�u�b�#Ξ��!
�8�4�����=#f�M��=/c>\��ɬ;!ʖ���ф�:��)�u�]������-�]}��T�%������YO�@�8��H�֏2:}:�i���m��`��k+N��]��\G����|8�Z�Fjʅ���d�҇���������e��+�Ew�:m�t��!���Jo=�
v
_����W�ǟTd��C~ݲ�.�B��P��')H��j�"�v=F��^�l��k��l��ДO��R�e"�K=itr�T*b� �t&v��R.Y:��A� ��6]h��W>%�����=�3?sO��_,�U&���y��rL���/�n5��t�8Y��eTX)����b��q���0 �
�����~�qW�a�A�i��+fn*�_`��.\�C�)a���!{�&{i$����F�<�-ɋ���(�Tp+ǘ'��r����n:�j�HO#0���6](���q����Fl �q_�C���OS&��Q1}QNIp���E�C�H�u��5E_`���K������`�ϲY@{8����.�L�Ǯ�)���5�i��Th,5�P�@N�2'hi���iծ�����K��z�����o��#��Y("��ɹ�3(� ���"-�U��m��d��:�'���t[�:���'���~�z�3A��a�!J��O�ØG�Y%��� �<���Di��]g�К ���۩��1BR��=WIV�s��t�N[�6/ʛ_���3��uDx��g���]!�F�t0i�����^B��g�]_�4����_oo]���Ԕ���>g�UN��˫F��K���ǂN���ݺ�ֵު��y�>D8����&�P礤�����L���v7��>h.�ު��J�K��$]Y���a~G�3��t��P��M��ݻ%�� �ea�s�&"f*$z��A�̢��S�!&�X�ajP��A�զє��?��y�]�v+ܰ��J�zk�h�2ݓ��^
��vK�tce�pC #�_z�1�������@��9wPi#��ݑ=��oZ{��3�|K�1�9PG��ƹ������3�\W?7/&���E]�?��B���z-@BH�;ʀ��H�iʥH��K��~�F��ׇ�4�����X9��H�?���I��t64:���o��߰|��q�$*maЉ�F�=���F�0E�_
��c��#����ּ�:�J��W*;�|����[��韽Y�7�n0V�Ѹ�#���
��ˣk��:_.~�3�HY�{���`>w^8�CG�V����fKx`��zmD�@8�2*�C�2���8 %Ps����
%�����ơ�����v��4h�x�o�$}~Yo�9��:3.u���#%��-�	%�_��#{�ﳵZ"x���[Q{�A��"�i�-�%AA���LK�6��u��2�>x��D9�:�d����m�G�=P�dO�C�,��8��$.��@�1������4{���,fzM�;���S؃������g]i`p�*Bu~uLv~�[�r�i>�*
�P�	d�j什0������_�@����۰��xSE�4 !���s�*C�Y%d�����h�F0�Nq�i�,��-�d�ܽ��94����xx ��+t߭�W��|��%�Ѷ��(J/���:h�$��̵�+Sh�s�_eb�[v�p7�aC��)b�9Db�4OEB��*!�Y0v��:���my������3|�J;`}��ɜ"9�o��OG9d�(]U�?g�bG���q7�D�+����R�*M�ܣJ&��2�7\�8wB�	=E���J��o�⿐� ��N�-t��c���D���#�R[�a�`�L-�0S�=x��,o��̂ ����+8yC,���A����ט��`�w ����IY��#�UJ	��:�n��sYÓ]6�+��E%�ͷӶ�)�(��G�ox�n��S�[��>i��*�Tڟo9�s���$<�7
��D�!\t�M�s0�6V}�I�VI�]M��~��̃��R���N(�cz�ڭOo?�ta�.w��2����g������jމ�b�T��]������SB����y��wC��m���.�AV�����3��,ASg�n#���pJR*�=W<[ ��4IU�D�����56_R�ZE"��%�%�
 ����I�CŚW�\[ݵ�\��7X�vzǮ��*�+u�4�o/UBS�`Q��ޞ\A$�GlMJ>�s�*F��0h7ǣKA�D\���Mک�2��������w���ټ�+Nťx�����j�,�Drۂ�I�}ZW�?��|Vm@�_��I?lMe/�g."��Z�&�z\;�9d�<(����F)��#��i�j5� H)P]��\��.�W
5k�AAX,�2o��
�x%���A���Y*1�_��=���P%_��Q_�oQ���lIa�>����d ]N���c$���[XT@��rF�3v.��0��Aێ�on�Kb׷���A�ߪ��w4��g��rd�ӉުQ���_[X۹��O,��:�/�=�a�����X�%�����y�6����6FI�衣�\���/h���f�̫�08]f�L�O�<d�A)q���R>[B��l������V����Qﵐ�,����y��I�+b@T�.?H@�r���X�}i��0��@�C�>��Ť:�f�J&R��~����VRXlxV65EB    d014    21b0��l}���`׻7u5c
�s̌Cx�:��+��$��O�@�5�%�0���<f@t��xM�����	Y2�x����lP�z�uTT%�O<��]�&�����h>�͐#�]2B�5`#NV$!��3��{������h��)w�����}K�����-�a��{n���1�C� �����4��yI�\��f�ì=\�����1b!R=�l�n/jpe<�2*�#u��R���Sj�s�=>�]]���i�n�X	9��EA��Ժ&k;B��y]����5}m�T��R�0Ǹ������&5�=�$���7�?w�7L�j��l�WW($,�L���Y0-?B`����^�)<_Mt�6�?6���p���rF��=��K)������ j���4[P�{*)�e/ˤ��q��!N��lڭ;�Ҥ�%+�xt��r�:3`Z�[��rI/���MI6�ov�pt��G�W �/H�OҺ��:1u�c2\Z���"�4i���X�},v�������(���侌�k���eM�����sF��2��d$C������䍼K)?j��(�,g��i�j�'��Ϻ�]7�\�-%��v�\�<� W��_m�I�fO��N�w9C1ܯ�����ܵ+m	#θ���(+8���aW�;����q�LpR�	���M�����=����C�+���p�u�V�1'Zz&-��A#a�vF��ܬ��Ԫs�����0�X����8�O�P����1M���p�.��/E|2qʻɴ��J�2qn2���I��Lt�ius��k%- #ұ�H���|2�rQz�JgA2���/�}���"?�Oz]�����(�#�ϏqJ�lf�,³=0V�jk1�?A��Y��I�>���B�����y�	�7g$+u��hZro���7[�/�1�j�1�L�<���
��,�]�{JK�,�~(��'������Y7�X�*����%�9P,tN��F~���c}r��IdO��'����E&�O		���)zT�����ib}!{&�˧�DҜ38�gS�ɸo� ��~p��"���"Q"��)6Y��������s���,���]e�~��y-d�iE��7�}�Vi�T�:����B�ӈ_��m�ߝ�G�z#u$��fH.���m��&���|�X!�����4)�`L�?�/�����<p��s�*8�x�܄�N�<B���G��Z�Q�D�����O`������%=������N���M��rGѼ�Z�j����ޭ$���uU����{O�*����U�N�ؚ�W�s��a�ʢ��#W�O���	8!9�!@�u�g��`f��ڝ��i
NO~!6D-�����S�s=D���G���@�pև�]\х]8�����*L�L�*'k>�|���.�N�Hg���E�X������i˪����*I<�L|ve��פ�b	�B�&�l)����7wF�ۊR"a91[�0� ��)�
ٺ�f+;�� ,E3{v'�xL����D\��������Ά��!,�(6�^ظ�����{f����Q����w\4�W�$<��捣txKc�E%��e{1��}�5~?4���4���Y�L˦����&�F]���{6U�Z � ͑�N$ba2��'r�8�%��I��9REG�}��2�{�'�f��$E�.�ʘn���!�5f�U����n�V����]\���=�DN���>�h22$s��qg����/UBnd�����M��z��`���!���UL8�56Y������Px��g;�o}���0���yx]�`��q��._���R&׎ݻ�+�wV�-��Y ����p��q�l���bůLP�w0l�a��a�2Du���E>38�c1�Ӊ�V(��:���ε|�?��ZvK��m��_I�1��z�����u���7(u���iV2��R.N��nn���Bz�����P���v�t��[�����p�/�@�k$����Z������+�nz@��ڙB�ԼcL��zy$<����|��.��8b�RG�4g��j$����FM�o;���'�U�S��{���E�B7��wo-&:���.{�p��Q5H�}t[�s%��||��}%Qz,�|Y1���U�Jr	Fت�S��UD��H���&���Cr��!��Ͷ9��L����j��Cռ0��=����^̇vA/��������B���,���U!|ÉC�t����������̇��o�ͩ��S��$do$�|���F`w/
��1O�}�~{j>�������AA>�Ozm���2�	^�\\��?���@�}��NX܊NS�:Hg�zh��u��W����AH�:�vX��3딾�a%-r����e���}]'v��V�>g�R���^b��2n4�2��bP��%�)B�W�*h�/����;f]����+ ��MD�6MNL���|:wN?��p'Hf ��"�/d�Pn{gs]+D#+{�Cn�WG �ƙ.��m�ZA��q������z�
��MXHٓ�N�I8��m���B�W�8mm���*� ����E,�>W��\'u��Z�ª�+`K�D�Rٻ�rJ+m�{��0\�	h'R�`��ʊS�k�c�7��ƲX�_�t��OsXx�Y#�#�d5���\n�*��o�D�îl}DWH��*��������B%*p�p~2A�����M��1��+�,�W���̭#'��5 �w߬�<R��a�������	��[Q���Vj:P{�K1m�C�����Z�e{V��铥�>"	�����Y�*�����E`��/�����b�&�ȡ�3�d�\yK����

P��=�� �N+Y�`���_��u9m+�M�ʫ�r�6E��v�뚟~F+�}B�	T�����٢�>�-S6�=�qE�)G�
M}BӰ��d�^Z�e�s���4j¦/�ҟ5d1YSM����@��M�����$=Jw~���SAJ;��X����&���w
DG�����q��!�qA�i�խ�_�f�$nS�l� .}H}CbG�6���7\�&�h,?�-�Qjٍ]���]c�d��@�%=Xp���(#lu�k��
�2E��j^�Jn�1��~�D�������mTO �����[\^֗jl7r�m7�$�$����,9���6"Ѽ�Z�jd9|��j0���kA�Lq�*�2�6����I(	�֥%��' �i�澒:%�CT���%l.��02�=���#��É�|�;�����D�%�z����Id�X�Ɍi�3�}�<mM�w+9����O�V���d  �Z>z��H�So�W?gZ<g��l֕?ո���@h@�wP
�8�v�9��a�)F�(���6ƫ��ȕ@J4��*����N��u�3�#h�x_����xF۩`s��YXd�Q,�� �"]�_ ����e�Gv>^7�K�#ݨ�?v2Ӄ݌͠H��p�d͔��_m��,ЖCȔH��T��< t���:~G1���	����)r�|_c"%j�\y�&����?%�ɻ~�@��L"]�,8Z��31a �&�Jb:����n����Y�HG<��5�՞a�S��ݷ��X�Lׄ��v��Pu���r�-�_�%>�>4����֌7g���g�`���i2	}�u�Et���,*��U -إ_){A��Թ�_?X^�U�ԣ%���Cy��8������5wog��#�FKu�I�1��y�zQёf���Z�H]{u��&�B%�� %��X^r{�M+V��T��'P���x���u����Ӳ�ϔ�}X�=�c�|tp<uA2w|���Da{�� ]-��_6���|�}���A�T�t�M�o8k�I�L�W�upBK��5NNP���2��򤂪	գ&;�	�����J/ �	�{S��HХ�]�B`�]����w�7��X5ͦ��J�d���@N�B涙m�4�pL`|G-"`�8a�T9��X�:�x�X[���(ռ7�(�f՘I�3[t&@2��
�L�=Ύ%&���3�|vP�����X�_WU,�"M�mp���paN�m�:W^c=��X>�m�l�{8_~8��F4��a��D�W�Z����µ������[��1�z����P�� ��+sA`ʗ�0���(OB��Y�N�b��� �5�K�v�x@�9�	���ʭ�R�R��8X��'�R�\��'K�:��ۋ|^�7�U<�Aһ���f�<���a��}/���B���C��Q�f�}j�#ˋ �{6/w�0كZ���V�����F��u�j�K�G��t��+�uGO��V��ן^������_�US}�	���
w.!��\hHq�,V]�$�����5Ǭx]1� �u���et��p�u���A��>-~��є����A�_�h����?�2)�Ց�?1��op�M#��~[�0��{5N�=�ϛ�������J��s̜}�!g�RW�X�%��?!�hB���
��	D����^�}s�NH�
������w1�+9 W�	�+�J��x��v��q���cJ���9`��@]ւ���t@?LW9J�䷟	�_@�k��y�d��T���_zO/H�����(��>�^"{wh�J���վVr ������|X��F���03��B��1�2��d���*gr�r�g���k�2搷����h�Eyt
�E�䴲$����e��apSo��\��Cfo�0��6�bT�_CH�H"ݻ
w����i��+�^�����N��J�����xP��|�d@/��V�,�DBi����z���#dx1}g��Z5®R��n��4@Ec��yC"�*� `��<����6���΀Q�M�Z� �o�G��� ���Z_�{AYG*)�=�޿���S=��%k���dg�#9����r�փ#�9%�FR����hX
K��}#y4�I��m�`�bf��h�eJU�AZ�UD��"��5�3�W�5H�y_J��u�n[��.� �g���U#1�{̔gS	�~�q��@��ʠ�C������v�&5/m $8Y1O�q�vͥh_��o����3�o�5���o��b����\z��h?FX�|�E�	c�e��4Ŝz�`��W�!�X]��k�.2����=����䂰Ȝ.�gx#��Cߪ��w�$�0�ʞq0ߡ�6�������
���jY�6��݈i���a�#'[w�5�"*��R'1��D�Qp����T�[I�~��˨ۢCHq�	>�h�bI|�m�'��٧z|��Ryr�9dc��$>�>��IG*�\����[�XӔ����4]c����1���祾�{>kO�>clc�֓
��%�9���A�n�;,���ر�S|���Yr}��aaj��N���1]�G���=�O�^�uo�-����մ�dK��l�b��B�
%�l�&�`�F�⪧lX��yn.K0��nf��y�LB��l��_�٦�l��S��L��7�� �L�2�g��1'��FN�J���&�O%)���}6W�}&�1,u��չ��ʭ�� �ުP�zI��F����v���2�"��n��<!Ƀ�lW^+��&ro󸀾 E��d{n�}��0�4Sʭ�2i�?ğ���[�D�d+�?l�*���`��4Ћt�+7L�a�r�\-y(J�*��#�d�Od���E	T��T6D�99�*�T뵑�� 2��VA���M�[6�H�^���'.��EC[K�iŢ$�S|֚��DEv�(���V´r�#Im�����]~�v5�Ű(�Ɯ�lS�� osɔ�^�<��{�>0S��&<BK�mD��g��b��ogVٷ���)��ʰ������MF�#�HE�"��% �+�Lo��{���٤$��<�j�P�f߮ߋ�jT]�@�.ֺ8���[o�%z��^��'����$vr��tu��&[�5>��{�)�Wy�~���c&&��N���:�ʚ�j�o�����a�j�M]�� ��P)d�\G�F;�!�'}Whk���s�R`EW�^�7�u��ו������.|M�R�)6����%��:S+k�rM����u�Y�f-�g@s⁀}����+����6F��oX�,�S���B�y���{_�v9v�}X�����H����)"���{���Q՚,�V3�d;y)�1'�>F��K/R�5���`NIk�~��~�tJ��G��7���q��6���_���:%���2NAY�\�.�g2p;���R�n�d�������!h�Z2�h�AH!B��b%T�P���}�e�G���xUx	;5� =����@��6(fS_v"��s�Wq0%<�|'�ܠl-�e]���\��1^l�ȋ��zE�},ݼz5ٺN�m̢�62��}�仒���>�ܻ�4W�����T"#z�Mm��r�㻀���1�|���w����	m���ؔ3QP�n�xV�v33�O-�;۷61�:N����8ڪFNڀ9�aQe	P+zxhЖ�ʋj�Gx���g��/�.D"��2�cX�'����%�EH��$���k�o�4+�3��B�ִ`�2�Ù3�P�&�XxJ����b9����1��L��;T������إ)��(�5���&z��U�BB���P" ��>��A"�h����s�D-�����O�
W������BLi��#ʍ��a�]a4����).`0���=�f�N�A�|"ǟ�t�� KL&M��=�#���Y'�YGv��9?�f�UW��?�=���̗3W٨o��8��
N`���rW�Ɓ����_)K���o��MA�-�:�H�C���1W5%p���	�ؘ������ь�U��R~Pf�1��uU�q$�<�0&Y �oA���K��� ��N�~�#6�Q(aBj�7�v�R[�Ւ�4W[�����x��|�V��X�O��W���ZԢ��֢���o�t�,$á�m)�f$]�iH%�pL`~�>�*H�R���Q�x���0��Oܓ}�^��O�r�?=Fnk��9��I��a��§�"��=�/dZ�oF9�v׌�E�}��v�>=&�~e���u)�f.��� ��Cf�΄�:�w-�>H{�X�<����N�Av%��_��5��f�'2�4�Y?���KCHG�̊_1�F
kQy,A�W�s�F��<^3V�6K�{wəG�%Q�//�Qm ]��UVA�U.>���,�W�.:�;�W[F����o�~��-�!�a�ϕ�wJ�)R��g��H7�A��2ư�I���k!���q͢�@b�8v����K-9��@�IN��� )g�xP^g�i{��������8 ������Ls�x������zwp����+�Z/g8/���8�$�	D��s�a?4ʌ�˄�GEV\ys���
H��fѣX�
/EO)1�S�8����f�A��"�a�P=)�����7�8�įT4�v�bcF���}1��9A���5?�5qt&�]�4���BBJV�"u�
A��d��^�X���ͳH�W�r�\3�R��s�=ޯ���꘮��&��j��:�]t9{���9gT���"��2Î��>ZF
�ND�}ys�&�=� 3Uk�/Լ������D��ԑś#N6��+����ǥ?A0S���O���]A&(�f)K�3wX���Bm?_�(�z9���S���pDP=�I����t�p/���*w�`��s`} B^���L�2m� �h��Ȝ<2Ύ`ٽ(��M*<�x� �=�n+m���A�;�͉k��p�~�J1������GI�!1R!Rf����j��Z~n��H_����jJ��J�M�Fʦ���'!X��;o'F���Xy�c0%�sO�lT��O�"��z�u��f��@Jyf�>/�5�]?�|����I��:�'|��mjL���a C|$Z�2!8�Q������������?�����+��#7^�6`��>�u�1� �M"�ơ���\@c�L\��ˀyk&�ݑJpo}��"5�#�Hء�0��k��c���z�#/�����U�4��*� a�E�brD�=��������?*�� .%e5h��`�&�u��G7�R��1s�������* =HR�#�(7-��39w�PKT��~ �2���L/ۄcZè��@i�:E�}��Ѥ`�ȍtb-�D���Ol�*�$]���o|d�j�/����~�W�[sE�MU_��,�ç��{4�;>Q^fk��<�	���e����R35[A�L�F�����L�\��I��D�@5��B9N��ӓ���=.H����E�.�su_M�����X���j�������N/�G��f('�Y׈�)��1Z�� �x`��mt�d���ÍU0羃c����Q�c�~�g(&ᢳ��nV�)g~�]9��݀���L5&�-ӷF�V�aV@<߰7t�����9�c��eRy|��yxZY�&(rSO��F�T�JR�g�X^o*!�Ǫ\��#���p]��e������2B(���T���,�,���a_U�
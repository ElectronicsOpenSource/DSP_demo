XlxV65EB    fa00    2920	��Wt�,�֖w�n�%�!�,�7��I�U����$i`c�  ;̊Z�Q_i�'^�{	����5�!��W�H�$� ��X�4v�L_����Go´��T|����h�J�(z�/���bS�ocVu����s�B%rA56V�(��rCD�M��).���{!������A����j����O:�~�^6����O�9E���V���j��Ru[1�rnPS��m�p���i��,ܳ�t]N���_l�9�$u�x
�_3bE\��GH.) ���_��N���B��I�FF���x>���E�$z�I����O�kl5W� ������(�OmK@��[�eG�b�Ȗ�)!�̅��.1�m��8�(a�s�ځy'EV��%y5������[F��x��
+�K�D��;�$�A��C(.MAb�N��'f��ա:{Ǳvzr��@�Q�¡}���*f����X��m!��ޅ�c���6�s��^i���O@U˄N����e{�g�VeR�jK��^�EA��h�oUt�-�r�Б�!��A�w'�0Ϩ��{3k�����Y�r3�[�z5��+�J��;�$c s=2&0��d>�|�TR�"�F;{��)�K����^z.J����^�Й�Jh����b0Z�*��G�u�?k[���*��]�fр���W  �o�s��+��@k�o�TF�RT�bu�ȳ5����Q%, *e!̦R�C;>��b����O
B���u3"}O�ʷ��"��Ф�����?> |��s���mt��i��V�u�q��E7�] #o8�H$RS�t��)7#�Yܫ���s����#���l��"?�&�[v�oƆO%�^��1�	�Dˍ�խkc��
/�����'[u[���݉��'ϧ��o���O��Ow4��d1D�L��=K���U�s�������h�f�����ثv�N[�A	9�m�r��5�oI������,��]��fY�'�?�!Mfn轿��+��*ie���կ��`��c�t�O���sK�����|�PJ��8���S����tH_�3d�g��g�Cn_�E����F��C�ˇ�U�АQ�r�!��'xZ�ӗ�\6Qy��n[.�eGS@��4Jh��Lܯ}F�f��k#�{��s�F�h)
�M$,��}������P��w 1π��xr�o&+���:��|k�Wlr�DB�b���[�'�F�	@��rHl��Ʊ��מ겱��Γ��PU��p�g0(�z�U�־AX�_�־0���+�w��/8�\���r��2T|�~�}�X\>��D`g�n�"7=��:��6؂M�@j���O	��K|Q�k���x0�x�V<�c�$��\�~[�"9��dc�+�[|����k��A���M��Ȳ�޽�f#�k�σGP]]�:�����X�����N��kdH�Q Wk�2jB���x��,Y��K_zg������D��Z{?~�T�s��_~�����ү�r�F��/�xҭgNs�!U���[�7Db��Y1nmN�H	���3���V��0{Cl�n�?7���2"ݬ��P�b̭n�^JM5��q�9ݥW:����8r� �]�p�6a���eUVȳ� ʥ|�O�0�:�ܠݾ2]/z������J��r��6�vx�/K�?r�o���A����Xઞv���Y�]@�^E�_���%N�
���(e-]ʩ���V�pi�~��VT U ��ĒwW�N�l>E�&g��̯.ilő{g�JW�R�c��������[R1"d�"���enZ�Q��՗��e�#|��ߟ^Q����P�r��-d&�|?}cLyS��A�T�V�W"������G�5h`�C�\���s����Fm6	��?'#M�̩A��{;Ü�����=^R*L��ؒ�f�"7�ڪ���\��� [�v����˾BEH�ʘw��P�*����י����JAq8a���2S�h����Ƒ��Ad�dH�w���:�	25-=�vb�<]�a����j�{����9��+#���jұ�����H!��@����3�U���v����r��Ԅ�}m�'�-��7����s>t��	���ϛJo�v.��k؋��7\���y��V��PT��?�Oφ\��G��/�wS0(3�ە݄�-�Q��)1 Ujvm��]h�%���}���ĳ�Tb��z��?�_�V�deXa�+e�r�Ӄ�n�TՋ�M,�]B2��-L��/K�ErTmuҰ%��-k��#p�jx�C����f�}���u��Ԅ���2l��]�>��N_��m�� _���s�,M�'�\-�����>�.�1�vi�t�� v��t�<�B%��J@��4��@�hUYk���-;�,>�v�a�yM������u`��VwrH�Hy���7�E���'x	�}_�ф��I�ȃ��mxL�VK:|H}J�N!��^��.>�7ﾮr�ZX��-	���XR�:�++y�
�	x�R�/+�d-C�g����7�B�^�uΏ�=yx�û�C�	*{5�'�n7 ������,��ڂp��.X����w�}��F��#q�����|�"x�yG�s%U���g��a �{��֪!����3z��r�4�4hx��f���pcβ�9�c�Ϋ�Q�n���_��cY}�#;�5º#n��E9	F��@RW�[�����bƝU����)-4v��tqY�By�mz��HX?��@��� /�^�5\��-K���g�����%�l�&)�n�ybŃ�bw?=�iO^
Wߘ����7(u�?�(��b����B)�ch�/���I�Ӛ�_a��cCl��#=��o�&�ؖy�Q�$�i.^�nU>S��@�r����N ��!��j��hAk�hnH��V�ʼ��*�Z=�tv�V���R��EG�Z!~�,53��.v5�}�8l�K�1_�9���<����ip�`7FcAt+%�׷4)�Q���Z��0yQI��̟գ�9W-{�K�� �*�0�z+D��9Dc��[H���mj'�߼�ҭ�qe=0,h�\o�I�	��?�g҈k	�h�-Bo� � ��W�`_�F�����vt��~IE7�����1�{#S{a>/z'�A����R�	����߲�n	�<���\�q�k<|0��sHr��| �h��SU��|㒩Lß�/'�o>�|�=�q#�;yI�p�E��ɠ���Q�Z�Q�w8�^������Haf~xI��y�ޑ<��Y������B�x�IL��J%A�q���@���(��>�W�
�=�܅9�v��+�stI�h_l�?�/��U�#�6x�&���ňG\�(,#��t��� E	]��Zml����YK;U!�m����j��	�/U��'����X���^��?���EB��q�5k������S���1%aΆ(nl1٘4�8��bv��a�$�:�*�����9|$sG�	w׎�ζ�r�K@/:)������K�O��Xt��O�lƟ�&����E��+�%+��܏%��E��_iz�d[/"��piU"�}��"�l�"A`�؅�[w���6F4�ja�6$B�jn~�ߞ�p6( ��+�a妛��^cÜ��l��o����fK�vD�Zk{�
�����Tv9e���'5��!7�<��5x���a6Z@E�$�Z��G"A2#)>���_sy�����w�x�����?]�t˴,j�&�B��e��J5���jx�.Gt��Om˘e�$T�	C��U�:��ԕNF�8Cuw�g4�bL�@l�2��[�	�# �L�E �W�V���	��'���FH`�)a��!N�1��k�crH������Qƹ�4Ɣ����qE���g��{j͎׼}W���.gÞ�F>�_��#���,d���6̥)�2]o���e���+˃Y,��3a}�W>�Z�S`_"1ixo�
Q �v�'P�� �<�t�}��A)����Aj`�N���͜�-�����"�^��
������M~]Ow,�a+ll�L�Z;��Ԅd��)ǽ�r�����f�J�R���r��+eF�bs�	>��2�	B�;k>|�5��D9��Y�Q&t�7#Iz���M�9Z��+_��r�/Ȗ�	���$T��\]P�g���j�?�������@2�wi;����S|������5^銙3j���*Q�z9�=JP���p�%=�W�fk�s[G�8;7�q��Eb(|0#]�� ��W*Yiɮ��N�w`�^k�h[}N��P�H�,����:M<H˴��!�X�Kd�Қ���-#��}\e(�QH�bZ5��e�.>W�.}۷o+I�;���h�=m|�����~^��!�L�vq�'�6%�O�$V|��a0 E�j3"��!2/�����G���ѯ=��mGP�R`A���p�)�V�ˀ��IS� .�`c#�Ї̄����㥜q�lh�`qJ���;�x������c��V�g�R�sy/�����CD���w���<V���k�`�I
�>X�B�x��=��V��O�ol�c�/e1��]�������ZȆ�I���Z�+�*D��� ް����9�PjМ��LrA�H��"a�e`�4���WQ :'tU�/K�G����2\#=g���L$�Y��tL�����aB@�yƈl����&�&Kv��6�{Z �7s �S�9$��Rw�Ya��(�`s!�k@;Bd/���� ⶉ%� �����*I�R��@'�a�&p�k�<�j��c���k���@�:V�)�Cr��X�AY-��[�aW�U!X`�P��=-~M^U§�g iQ��ϐ�(d���TqGx�n��'V����S�6�B׫%��B'�����r��4���]Z?������]��]''g��gzĿ$;�����5�˜n�Ҟhb�	]���^n�e��hw�U����0W�"D�G�S�9�zh�D�=��L瑾)tz{�ԝb3�G|�@*,�T��y�� m��ۛ^hI�_�c&�K����`�=<-�i�n��~��� n��D����ڡsփB�נ8�-�ٱ�)��>�ޜ���<Il�؃���'��v�r^k��wZ�F�^���[����<+ㄙ�����W��ˊ�Y�ĩw��_�(�W��p`!���5-'���M��.�	-�,㕃*	f~͛���Q�v�D
�Aa͹�T���_Ӑ�*�me�R��<��Wq���h	�dm ��o�&���B��۸��Ϣ��c-��U^�a�J��� ��`'��T����l������ԁ��]E�d}" ��~- rwIυ#v��%�Zd�ڇ9���ӵʞ�}U��)�1I�����H-7�d�y��U6�)�\=29v$���bk���k���1��7*_b� Ϳ ��]/�U�zo�t�ҋi]��k���������<g���J������܂�`8!F{7mфj��⃵ܡ_���Q��$ٺ����p�hή���v�ju�=�/�?����;:Oz�(� L�w����;Hȇ����)�c'��~�p�%��{&o??cv�A�/�/�a�%�e�=��L�������EW��&��Y��<cM�)�85�� �ùu�/��s������\
t�^�������z�F��̶�Ѩ(_�>��ʞ�W�CJj��'2懧�Y���K�0.����|l����O��H'bL�@���O���V��7��P���{ݻ+y�M�ռ#F+�;8����z���d���4U�A/�te��!�>ȓ��|�OPY?Qԧ�|k�7/ �q�1la߾�[��n;�9��A4�1�Os[C����ݜkC�cqJKg��v8���m_2� ������*���P}��1@�[qhte�$�$c�8�W8��v�y�z�"MD��TOT��έ�>�mh��,�He��,�Bq5.Js�?H:�qT��9*��e���?���������̖%�t��oEj��R	
���=��~��#�O��/z$��^�_Ud���==i_���T�&յ"��s���u�͈�!H�z��K�dB�jhk��K,d7@Q���&�|s�#&�w��/����f�fB`�H�OЏі� ,����#�i��N�(�3�jm��M���<[��� �Bk�8,Y; -X�R�X�~���Pwj~Ӊ�Vfs;�p����"�:������!l~)q�T�a�v �p�o:x��I���S�wg2�f�Թ��LcID�3���4o]���K~[��}�dҺ�(Z9!��VG�bEؔ^v�)����`5>D�Z"Ű!���z��G����*T��ا�"�t6��wpٞF����?]a���I Xe3Q���陰�\�}P|ܲgb��Դ��4��G\�k��ݨh�:0S��O�T�v�?���U�9M�����z���Ŀx�R@��<�if[Ȯ�p�Ťg���g��)�����VwI=��R����(�9s�h{��ӤdH � NO�ܵzI�ɔc�s�yb'��Ws��c�]Ψp�p
N�M2�j�J��Z��Ӹ!tu��'�M���`�P"���5 ��X9Ե̟�'�w�4[��Y��rK�]��A�b��棷�T��=�D9m�g(`��o�
xR��*���EX!US`{O*�ꔿ�ړu����*����w�B��v�E6�X�� \$Ϙ��q:&�_L]oN^�Yq���e�5�\��s��]�I����n����U�~�o/L�|ti&��L�+ȍ� �F�D�7��I>z{X���N'�<2�w��l��P$1vO�[3vg������kO1x���A��Q����h��n�&M��҄�>���ըb1h8�T �΄@��T��BM�#�� j���!��`[�~�N�;~Z�M�<��9�����Oܓ8���it�\��=o��N����;횪)v�8��T��!w�0w�j�O�bÇZ
F,�`Tf�/�s�vF=:5��nT��@��g��ғO���F8�N��蔙S�>�p��=X������-��>O�0R���Es�h�dB<��V	������ȍ���N2N�+���>�2�G�E�c���z�G����E�g�섷��=y�n^��u�$w����[�U�_}2�m��YP���[4�W���0�����g!�X�bδ�FT������E�sDϳ�o�Z�b��0n>i���7�+T]�;�uC��߅�n��Q�����o@�V�&�����x�H�ydO*�T3�o�w�B�Fmj��1��5A���*a��t�5C�
�|^�f�ל~�����]�Vջ��f�c��,�qñ`����Nd�������w#t�O�b�˔�"a8�cgXR�2�AM.U8H�Y��!�L`�x<���rNٯ��D}��#I=8[ 6���wI��� 7r���s�02�]�W���U�r��������&͗�:��I-��"^*�����YCF9��
8���$e�C�����L$`��)�_$&WFA��JN���;����H��]�����U�d�u����fH�jߐ%M�N�u1!�G�Q�o��3ƲI�~FJ4����-�T��V ��K{�o������R�垑q��u�9�l�'I��)���K/�΍��0|W�Kyb����c0��4\��R��aƕͳJ�g�&^ �%LK�O�E�����Uө���fzMc��(�(�(Ba!q�ⱙ��0#\��Pƙ��q�sq�RM��6��,g2���o����������R��\K���,�7�0�K�f����Y�x���gA�K\�e4Ό�nq2��y������W=��݅�(J�p�&���*��F���
D�� �X���]���ә������Y�6���P�yۄ�z���1V�\?㽖�M"z�\�}��l~����M�͸����~fG�m0���sD����6�71�� ��"�,�u�2�
���׍�-4���s䟞+=_CoU ����s׽�3��w�u��z-$z�q�d�6�c�ODa�תq�
�����������8�A�&����&�Y^�������f��Vr(:��V����5ި��?����O��^9�,�vRA�uK������E(٭�p_�k��zE󿍳l�亂a��R�2�՞�̪�@'"�b�&�j�QtM���S�cϏ�D���hmӶ*K>�j�wF���W�f�1��N��扻����O��f��PW�$�G��fOU �oۙ�g[5���m��m�=�����>��ߚEE"��\ UG
!�g7����0�n�ků�G��6�Y��{��|"0�u�F�����z���UsA��'O�h��1�XPK$�Ȩq�O�����T[��e���]b�~h����>��_^�^�62��'sF�B���
=�-6+��Y2cׯ����ʱ�'~f�A�mS��Y��
]�F���qͣ��?�/�&ع�ǡ��:9��H�Kf���x�e��8h����K
���;�\��-$����Q5A�O�`�m?����~���%�Ң4�Z����W��	��h��}��>�1�Md���`
��9P�xc/yuI��N�<��5�1��r�Mx�G8RoFE�:B�����C�w��٩rT*������|~��N�D����|WO_:�1Rs0�{��Ї�8�e�� �@�(H�>*T�xOM��)A�N�'��=jpj}۴�8`�pl�(�'�a@kmF}��g~[���_��|��'W؞3��a8����� 
������U4Fl؃C9
H����윫��<�>���iFs=b��w�fI����5��oB
;=G��B���M��?�]ώh�wF�S�jI����+\qgW���^��q�ڰ��z� ��Ӿ��� �*�E���V�)�c{�}�������5��&N[ڏ�՚A/��:��u�U+���5$E��������Õ��yN�í��H�7�]���J�z���H>�W��qB�"�EY?
�3��|TAr��'�mfً2k>��`��p��}�9*�ʎ�y�P>�Gw#V�_�X�T%�S��!&Du@�|&�������g-GZ D�,tebwufzf�pKg�w���i�1��!����J���Z� PwA�����_E�E�a��1K��[3x�/�>�YV~����M��+K}�<���,�k��8 ���@�S�/:�CƬpiP�ٿ
tm5@����J�B|ѹ�������Ӕa�ph�h��om���&w��t�ǟ�V�K]�?X��_-:�Cg����Z�ۄ��y�6$���3.�!@L��ϓ�ȼ76\Ɔ9q͚F��],���]���7�iÏ��\�g�}��P;AJ�*�ݿ��	�	��0XUӘ��np80x�@E��7#4_�NdA��r9����RC�̫�"����9b��˷J�KR.~b���Ѭ���������x'��<׷`������R�]�)���i��3{&1�?^�+�����V��c��.b`B��cR����r�?�lm����;�XMau�E��x�O�v�t2 z��I���ҝ���,���d�h��aH�v39���h2����=������r}����;%ŕǹ��zVH�s>i�u-�%�y�8	7�Oz�4>�M��!V[=b�CS& �U�r�47�MZ6=)$�!�HF���\o������l�?�%�g��o�V�
>���4��/z�z����+��KT �S��1@��b�*�D�I���yO�#���� ��[�Tf�f�ΰl=��~﫞(�`
�M�[���Bn?�@��w����Y���:�Jm�8�F)9!V���//P#��"�/��[0gM�w��0M��I���0����D�%�ly6擾<�X�}���b��O��uŻî��PR�)=��Qj�CB�=�[�6̝�h�q73��p7R%-+�����7}��r7����GH��K��Nf���i��w��)g�r?Ώ�t����ŤK��V�85�	�����*ox�N����!�q߈BQap�ߗ��*���r�)�����kd�;��~��kxBO8
��8Z+s	��Uhh�l�B��R(�����h?W��2�5�+;��fN����<�mI�nSD�oWC��"r;����1$�;�Ɓ��f
�^���~GT�j)��/r;���{E$O�<;ên���.R8�D�W,������G��CH��"��j�P��m�
�W-�C;�o���V�ܭ��h�va +��PU�gG�G<K��L�r�ꟽ�҈w�4�_⳴3�R�����ޙ�j����Ě	'gL���s�Z$.�#AN.R)C�u������;����� ��R8O�XlxV65EB    1e73     630������"�K�*$%m<�!N�-�e'+��-
y��6��Z�F<�K²�lb���G"!a�i�5��;F��Ej�P�	�@N	���q��^T�5���J�ex��  W�p!���|���
� �-.���t�W-���m�i_�~3�����B��$Ɓ�D�9��Ʉ���!�����y�pl\w6O���J~򧂁:�G
�5$m�F��=-[�:s�L��:b�VC7z��n���*#��k��5����Ɍ��Kl��l/�H�,�#�����"��h��A��
�4Ǚ�mթ���YΫѴ"c>;"e����\�Ϡo��2����~�:��&\Y|�I`b{?�y|PT�Gv#D�L�H`܈�#$2Ѣ���H.(��~8I][��ݠ�bT�P��%�͂oe�G�ƭ%�3������ B�BfPug��}�ON��#�8z�A���j���0ZH��Ŀ*z�aϵUb"6sصlSJ��]�*X-��*݂�9n�m��VϪ,�78;c�)����ɝ;��kn%�(�������1Cʓ�w�$�Z�Y��<We��fgC��YI����?�B��� �0TE�Ȇ��;ϸ}�����^iWql�9A���a@��)�Z�[�NҜ��]5��'�o�����4u9�{M�<��py'�ЯD�ɀ�;�f�o",���#�\��x@���3L��b�'L�f���бZxuQ�� ?LV=$�6�3{�G.ls��>1ab���<b;�%��JA�j��Ld~G�E)!fQ'��$�Fy&k<��Rߡ���[�B��[���OMｌ��I蠟k�DA�h,OΩ'g���_0�N�Q�N;�h�����aE3Y�?䈀�4��H�^�FQ�7%� ��N��n�ӎ_'7h�1�7d �:2�9�=Ʌ��>��by�buͰ
P��~t��� ߃��Вp� ɓ�^�n<���"����:�iQ"����� �Fc!���E��#�����w%%x:��<ؘo+&���Y��	r���?=���F�{�9t 4���'���E39w����dKS�3O��Ҋ�I�5�V'���xF�P��Z^\9D���gw=��{�<�q0�:㚂(:I���=�Zg@p��y�
��=끩a��CJ�F�"�������\����'ś����j H?Z��T�0�褶 %�m�磟2B�����]�1wKFC5��7�3/����Q�H0�M��Ķ�e�=����e�����&Wh}MUT���lIt�n��$�T��͒��ֳo����G����!�������i]+!�P�����|������s:'+b�I5��������������x�ʔө�3��?�u3�H��e�y������S� ��<����L��.��ٟ^MW�Ur.�2�E��`XIG�� ���+�4v2�LO^��;@�Z9�5��T4+E]|��4$[��M_��ϼO})�Cn��;��$+,��T8��P?v8/�/XHt3����?��	_P\��v�f��6���P˨�}�VB�ݗ�����a����h�I���[�Fbrn�F��e0qY�����q����0��
XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����>�ߪ�ԗL�������]�˞tt^���k7���"��AK�p.4��V���1O�'9"�jEa��`��Q�>�X`_88v�?�%_p��r��[�!���y�AC�hh䡀BhQ	�〓{Ќ����W�)�H;vay�^���t��J�}��0ؓ�"ղ^)$�"<�����`򐠓�jRn�x���i�P[Z�5,[�Ј C_Z�T��@�W�d�� r�Z���VWYˡ�8���Ft^��:�K�M� �z��H�ڎ0s�����TuYʝ���0F��:A��i<�ד�I���.yΗ�S��9�M���������=��P�`�+�N[�h\u#e�SGAf�L�����DH���E��ʙՠ���l�3]���c\3���?-!�,{kMWc'��Z����)f���V�r|���v�sD�o�}ʙ�o�Ow��N�*Ru����e��L��	3����iZ�u�»>f�2���g��ģ�ۇ�2��=%��n��|�jyv�0�r9i���}W�_I?cV�f��T��d��z�/�� �%�?6��B�y���������҉��;�~�6p�����H���Ce��X�Ut+<79�,&��
�����F�y�D��~m"2�R��tY�7���D�R�L�D2�1�����#g�B(���f#6�L��H��%���,����i��b����0�]�T���^<�͍��7����@�)��z�ьul:�����q����;���XlxVHYEB    fa00    30f0�$Le�A�l��7p`�	�Q��z�P	i0E�9Xbc)A$�2��C"��ea'�"� ;���Y�ĭ�0�L~�����;�u(<-�N[X�*L��o�3�
�5�2����M�u���͈��k�>�Q/\�0�����N}&+��s�R��|՝����n�K�%�-9F�޺DR~i���+F�])�1^���ȁ����-�(��w�:�4k��Ok�I�c�����Y�,
s�}9^\�Y���}�.�^H�Ih#<�!Nф�]�c��S��'UNu�&}e��M� �B=7�p� r'��tLKm&G�C	��0��mM��y~� t�}r_���Q[����G�v��7k�©��jN�r~$�[ő�,[����Ξ=�;]�>�b��������z|�-_(*�ƍ�F��?���okB�ou%T�����ۮ'���ZG���nO昖 ��Ө��ry�g��r�v���z������Z,�
�dm}K��V�B���,{E�yܖv������z]����[gJ������^��}i��|�$�rF�M9|t���.�l�����87����0�y{��e%5��<a^8�#����2R��>��&�'X=���ͫkb`��b�Ӡm^N��θ?�͘`��M�Qu�)�{�#��>"�>�6���9����������\E>?#�ˊ	�x��������i�V@�`��O�1���������m�]uh�H�E�5�s��!��WC7Q�������q�ڀ��ձ�R8�~�o.C�|��O"�4����D�����̢#�%��%�pfsb� ǝ�h�6��k�K#��]�CA����� �e�a�w�WEj`q����N��=��Ŷ�F�R*�C�L����Hz�䖽�D7O�&�4g�)"Cqg�E�Vn�jpkT�r(�����
��p�/1	ˁ����=˝�v��a�+D�lOf�_�)�Tɻܚ������ƞ=�ml��\�i
�zjZ�>R��YM:�	��.e�M�y]6��tn� X��"���jS񨳰d�Ʌ�?��I0#��f$ɛ�t=9�Ҩ�.Ѻ��Uz�7��	Y�Ù×q��B�߸Μ侷|.82꣑,�/���͔������x����j���(R�r���Y�]�|M��\y������E�($jT��؊�����F������#����^9�
|�t,LL�Z�~x/��d1�m�e*�(t��e���L<%��qj��{2�.I&n���D��Q���?k>,��b=�_/�P��;=W�X�)����|5�%K���ϲTD�F1�Q��J���2�1��x�"S�zZ�Ǻ�͌�=-����*��J��2�A5*���֐�1ፅ����^��S�B� U(�������|���?/	��ޛL3
/Tc�x�MCx��B9P�dI$�TV*S��UK�K�ꆐ��k��5����-���e���yv�����B:���Z�3P!������,m�J�����Ml���"�qY�\�S�w#��vs;��-��J\����~�֗V)oKd�yk�aǐ�Z�̥5ͺ��5`��"�B� ����
����9����D��=f�	ׅ�����l�X�1_�ƆeIќ�f����َ��GB�L�G$ث��q��H��g3Ol�����wV��au���w��:�WR�ň��2ц}\�C�fo��ipղ����1������9qY��@0�s໭�
���p��=0��ޱ摜��u(k_
�w!��-�:#9���F;���-`���D���v�Msk��	BL���m87n�_��{����(��$�&�8.Ѡ�������o�r���9�H�,-�����q�\��?'�:�^��·p��zL�£R��p�m6
��d�{wkè���!:��]y�V�fk�Y��V��aSJl&k����q��암���h�+r-~����}�w������ŔE��}b����3Hy�I|5���}ᤤ�o&��aR��0�+�wf�ݱaH�4�>�����.Q�X��� ����*�ɞ"������b�Q��|��s#�]%�끒���ǯ 1]��'�t�v���V�ӗh�ncL��
�)�������ؗyu�C�j��Ċ���⣦��]S���u
$��ũq�
PȖ����g)�����T`������R�k�Ѻ@z���.S��g�b�k"&��n���}�z��x��G�J���{=9*��6����$�ޚ "���!k�����q��!v�����I��Ug�"da�W>m�w��8���!��~�.ց�I=j����
� 4���rc�ɘ�]���*`N�biU1�H���/eSKw�Y~_:��ʬ?�xo�{�^�M��VKY�0֤I��%����<�y������j����P4�jd��K̙b��}@@#�]�
J��6�J´�6
e�\<�"7M�u��W즁l�o�/�q�h7���ٿ���@f���KM6j�w����ck�CQ<�'��譓y_B�I�y�=1��O�Q�YױP��cc���|�����;ֱX <Z�������&�P�f)�>+7r�y/]Z'�d���,y<�9T.K�)G�!�E]O�����1į Q�C EF����n�qG�����:�Q8)�~�����7�)���2�?}ӘP��y�.ڻ=��:����U�ʀ1
�� ���ɞD���u��x$cq ��3L�Ѻ`��H��l)��s��
��������Th�[D���# i�X�++���&�z)��m�v�k��m���[��%-�%�F����M�9�+˶�o䆃����E.7��'6�����l�LJW���Y��"����{V�^��<���<9�a�{��mW� <�]��G�O�⃤otMA�5������=��+��N�5�8ʡ�}�S�,�z�L壝�M���8!4n��pJ\d�|��]�>�7�Bj��\'�]�yNU 0����9k���T�m���?�n[]������P}���J3c-�3�Vp�[�Y��Ѥ+��A�s(�4��({c��Y���Ws]��x�a݂�1#�:W6 C8E�$;-�d����)\^^�x��g+������ww�m���k'ܬ��N���ݓ�Y�%���d��gC_
-|��?jW��e�݆(R��T|��k�n>3��%��m��-�P\.	�2F��jӨy�/�q���Y��}����5hg\�٠�]h��]*��H�Pd�T�Q�������L���m۲z���.M���#�ؚ)İ������sDsq|p�	O�(���v�[��G���B�Dl�f���+��o{�������w�gm�KS��c�ضHU<-����δ��Q���l��o�s�e��u7����dƥhz����Y��۬q4H�$[�.���NՒ���÷�h��5VI��|���mM�>�,�"�n��O��[��l�)4��g�)���|'�o�ʄ�^V�*y�qA�7�'D���#���|,�,�w��N��CW��&R��k��ĵ��+��X^2dx~��2��6q	҂�>w��p]w�k�Z�\��� YzTr�5a�A�RGZتm�H�@�/B	{ ��2�jAڊ�ڕk����S��\�g�1��a=�| Q�?�\b:��=�"8�����h���ϫZ?O�n����^��4:��C���ʾ`�pկ7�E #E����*x���~�P�w���K�KB�������Z�|Xڔ\ԥ~��έ֫���/�Q̔|g1�PC��'�
�d0�	zA�W��K�؜U��k27|sy�r$j,�	t�e�]�T��k?��ak�9�;�ؚ_��F�V��	���Z\߈͛�0��9$,]��S%A�������{��So��%�����$��ʻ�}�l�������Q�~X��J����x ȧt�����x�sU�2�P!�yRJMC�b�C�Z]x�ݸ��Rl���N����d2�@��*�Q�9n�ݰ"���Tܚ<}?&7 ����&������D�e�3LJK�ț^��y邴��'�}��.ai&3w#g?�f��{�Y�6��؄�h�R��k��(�|:���P�^p,�9IojZ�^�@Y80���	��b�1FY�)6	�r�[�`�2l����A7�gگ����c`y�H���Cř-��d��z�b���� �9��a�*iSqo�Ԋ;�/����n�!�Ė�	����u��g�[�jIyRG�@Q�-6޺�ΐ��m�%�E����̕S��Щ1#�I�Ǒa���N�XkD0$���<2�ɦt�q�����_�_g{�ܲ��X�W'��r?2rY�ȷ�_��z���g�]=XS/��dv�O6|��
<�&�p���(솁�;��`��Z�g�4�|�~��{��(ϧ������sfa�a�j��;v�@�~�?;f/U�]dԤCl�}��G�����c4 2��V�Rˡ' ����Jk����T�x�G�/����ϩ����d�<����v�hċ5k�:pi{�-�w�Ȳ�;nFN��P�.�WZ{S\O�k�Yy�������m;Dw{�{T�Ԟ�M���,�P9��ϓ��Ƞ� ƧR��,ծ�� �:9�����Hm�q���؎u��ˮ�gϷ׳�mgadKM�c�ttz�Ú�6��r=Ֆ[?}�i�՘��oZB��,�E��2���FSа򺁣J���
�������Z紧�M��v����5<	�<Ή�W�5-���z?x"�HCt��_lݚ�ݻ���������W�y�"��30�<�Ԥ�l�2^=��(�E\_Pp��_�������.��[ �Z/�f�YK�$�YߟY�v�܄��f<G�7�H���<���U�������#���Y�f��u�cH���nf�'ɿ9z̎n�K(Q�"o��Vk?�^�H�M�(
�>ښ['�T�?:��r�KE�k9�ռ�Y�TB�\���η����K*@:��?���Ҏ9t�/Nqb�R�:'�W�&%ךr~���\i
�����#} ��V�M�@>T�s�0�1 ���#�]e�D�i���!��$��~Fi�3����M�=`�*͟�ޝkT� wm[o5�缠.~gT�]0!��uS�M�E��"Q�
䢬a,��;������{��������&V0G��@�Ag>�v̀�gF:���eiC�`6�K����8��j(�i�����Ϗ�����Jn�Ĕe�n*u��{��5wq)�ǦY`���J�e�+�
v��\���kMq��@�u��]b\QE��&�+�M���}��k����'��V Ü;Tܭ�dcu��*�>�2��o���C2S�o^�S>Z�W��X��IHS���8�H[����;)����0��#s�[9�2E��:N$��m����ޞ>8M;�K'���� �
���)�lr�T���v䛟�q������B�󄫪=ߴ�+L�׎��n2�g�07�L�jt���U�cµv�t�ˤ��,�ɧ_�Y\��;���䤡�|���ᆖx�&^���;@�'��6�����{n*�a���Wi�lݪ�<�!�[���GШY+�׊m�À������X���lJ�xgu+���u@�Z�d�V��T@`�T�񬭐;�V��"�EBV�5�������l�կ������9maW����,�Ӷ;��f��Q���� >X��N@�v�mx� q��<~r��W�-8��R����Ā�p��[�����~0��15���3���Т;�
	�����-�0&�}i������Rk�LT1����V � �Ø�EgMv�M�*<	=\<��s]��J�a�7�B,ى�A�5(�"j�D�:��S���t��kdf uRww��!�ST��P�:���Y'���7�w/��{cx?��g���7�3+��3���]�s_k�a�R�}h���/͖;�@f�dq�U&*�sKeI��=�E������frρ��c/������;��S��^7zQ� �:o�m�7	과}uv�o�_=A��I~�6T��*I+dtT���	ⰵ�Z�ڪ���R�� ?�f9J&�ǐ%�K
��J��'�r�E8a".�zӬ(}�ؑ��Q��d����"0!̀^\��/3��gi����C.�ZD�J��� ΢�靖�Ƙq�I��7�g���+Q�%��%��c�;�?~c@!n�/_wM�ps���8��p��w5r v�*�'�6MU��ӗ��LU�y?��P���gf"W��D�e�nPM��b�x��jv�a��66��I}1H0|�xCY���[ix���&��cd��h#2�x��99�����/�m���13��y�������B���I�q�2� /�a�v=l�纡��<�Ԩ(��E mV��Z(�#/�]!(D�l��o��{#H��z�bM�?��6��.���d�JX����=v�.����D����צ�e�C8��&�Cll|�SFb��"9hQK�'9���
�/�x���2��x��������#k����,�W\ۗR ��Y�ȱi7�Y��+�ސ�_� 
�q/w�#2S��L��4��=�>�Pw�qi��fV>W���0"�?��h�f� �Սн0I�����W�/(X�e �}J�SRQ����M�{��A�q�'#R����"��߉l����lLɀ��
b�b&iy��j����ϒ�.�i]؃�"J�.5�J�B�;��"z�G�"���
�j���0���(bs�F#��¹ѯ.�q�Y,����!��"3c��$arp��َm/���>�������W2�~ү������.QLL?wd�V"5�P��|f��5�`W�%��$J2%��Q/��731m�`L�1H1�X\��̣{���gt�2���Qi���J�i�EQX�	��R�M"!�-v�2�a8��w������-,�9ɷ��A��*�2�$�.�L���5Rx)���\�X(d{�?��`����*,zd�1�D�һ9��QS�@p�b�|yvi9����J��b���{�8%΄��z2_ǝ�N$4��k��^S�s3�
����]M����zR���@+��T�MW���8�(yߢ*�-w���I>�4��)�
��x̞5�Z�l��VF�ߠ�Gha�������\JG�C��Z��Q��nGt�`���@*���r	�P��5��eҘŕ�A����zBq!��CN���Z$�}�0��g�^5;0�kI�-�v6/ӡ ���̺��Ϊ�1f��S��3�>)b�
��j��mdM�˪��@��A�w��ݞ��J(h��D�БH`cP�Z��	C�:|�佤���Q���y��9�d��r��Wю<^e�"��j
���/���~�|o_aX�ݪ���X��s���Ю"�'�L�~G����Ǣ�w��y�����@tL
&��é[�̮�(c��Q=��]�N$��eY`l�XWk��n`pZo���D�U�>O��T�>%��؉����K�h��wz�^��(]�F��Cl,�vmdQt�㔟��d ��|KUP�M#$[����6;(y���q���KT�uU��5X1H�s�`�6?\o�_��0+a��ߊ��4��)#FW�s��}�P!���� �����0�:��C�G�n�>�J��)Σ��UU� �g�́�p�B�4W%59���t�q��a��d�l���hF��i.�n��ҕxt� �/?l&�s��;;)fEI�`�fD��x��G��aS0�4�`�� 
�Դ,�U���U����*B��7�Ԙy�ZPbU�AkY�m�W[��o"C���"���r�2h�S�3R7�2ې͂:ӛn�Ӕ�����!��#�#$��I6&􍒰��7T.�J�n�y����޿%�!�ɴ�G� ��J9!���I�1�ى�{��g#(�	�cn)�9$v�-�P%>��k�^��D��4㫆6
)YW��I��#��X���⑭��ގ�
ӓ�S�� \��U���wI��ɵ���y���"616dג�ݦ��\�fC�����U�n�Nd�����G��Qί�ֈ��Q�(f�󣛼~-ca]��⫕|��:w��+�j�7�1ǳl��!�H�u����Ñ�n߿P��,��N4u� �,�:]Q��Đ�2ӡu���fK����=����OP?����꿽ed��;Q�ݳO����F���{�1�t9�{)Ty�Uv��u���9�H��m��(��r
�f�~���-P���[~�;z��~|
-1\J'(�˘[�eC�*��.}�]CU�ӌ�f��CSLgL�o�j���b0���&D�WJ7��P�Gӏ�pJ��a��K���^��H)��ċ�W���I%��Kz�����~�Q�{��s9錱~�ޔ��ه�LW�~�vc~�ݔ�J>�c*O=�:(�CΚ�� �]�{�T��ɝ��=�D����֗?��u���o��<����MU�U��9&��������6�繙:H�\�h7iW���v1�B�*����ٴdn�	��9ֲ@�-��FT�x��O���9ǔ�s��qs�����Y3t�/�G�S��u�aT�9�h�*�A�2/؛�(I_�ڙ)�?����2�C@@��ǴO�&��� *rxÔ�Ʌ��ɮ��1{�ɕ!���{���|p��f���,�	h?��
⯜m�~����[���pO±��mYXa��`*�U%FxrC��P4��©4���^s��O	bxN��+>cNF�m����^kד��5��.rtI�32]a��a�.�׃������	?�a��� [�U\�֏��l{xg�x���H��D���bq�����D9!��O8Tng�&�J?��Fqb=��y��ϡ�`���Z!}�p�������T2�B�&���^+hڪow��B~�!��Y`�� �� o�!���*�5����l���jsVCE��y���C�h*+�;dj���3S[�Hc�(s�C�^�6�X�c���tb�@)N���X W/'U�,����^�x�O��'�e�&4�;Ad�n�R�HS��&�a�`�)A��j�"^ː8͗^eJ}8�=��ԽS!&NM��8��Ǫ��r?�@"��Y���J�ޣC]��[	�1�Y����I��T�%B�m����n�YePe�w�����Ni���Ō=AB5�g���*��>�9�&b��m"p����c����o�;gp�u�o\�����*e��:����ͧT"��Y	���g��jr�4�R��e@����J �H|���?���<_��[@pۯv�a�N\��� ��&3ϛx%3[�o�@�rM��Ȑw�|9�nƴ��9��*��@g�[F̣^�^�����B�>~����l�q�H;��l��橶��se�QI�$a�^�.s��.=8$
�#��}C<o������_|I���Ob�|Qux6�t(����	M^���"~χ��>!$Z�����b�8e|
_vdA����|!̪X5P��b�{}L�8%���]��;����k���aq�$X,d�X\�\,�U��<��Qu���S�a���--e�U�ԕ-�'o�nV��t��/��D__�-#0z1��돿�3PIf'����!,�zC����>ą����0Δa�Ĺ �:\�J\�Eȇ**��:4X��F@ᄛDb�'ڹ��奷v��9^D�.�K_Rno���.��,i!����Ҏ�}?�G~���h������J�ŹP<�hahGD��c�$2~�rׁ��S(v�Ǡ̤p2'�f�!��4�f�@巋�b��2�KE9���2H�!�15������`
Zb��Wz�[�7�bRw�4C���k��ј�Ft�����gpt�T�q���"O��,S۟���a �3�t�!R�`��D�O��xro�'����9G�����{�ͺú�"̦K�4��aI��L���J�N��G�q�$���3�&�$LG�O R|� ��k�,�Pw���K0�B�<b	U�Hc��.����������V�E�����&�m%�t}�B�ʷ�-�'l2��;������Z�~~?�Od�H�x:;�tH{��8��"��S��	��ӂ��/�������r�T�6�c��d�a�G=�CԶ]>� ��b�=���C��n=F��Һ�ω̮���Wz<L~<��M�٣��lf��_A4*�;v����+�ѿt�n�՜3-��wCC�2$�4+Y*_��6�<��5@�E�pQ���J$+�rt*?��X���e��^r��u���
�=���$�S4h��@:��V�������� �,D�:�ù}����^+�{�/�|U�sg %b&�$�񥳄�a������<�H�c��FwE9\N2*�.�ㄒ]�2���h�K�%_����1C���o�R9�1�����8=�x��32���^e��J[1��bk\�%�1n���ʌJ�[�)���Y˵Xe�*$߲
��a5a��vI[�_����ᔝ}^��qr��U�4E��_2��6�5��|kVi�A�Vfz
��rvq��f;y6V��Gv=�D��J�f ������
X�3������}�r��s�:$�P��>����|����ձ�F�J���b���%fB�.�i��
������qN�d�"�u;�-`PC�x��[��$⹾��X`�v!�S@�����yIO
���c�0!��C�2�͔����[��	��4� }�kO������m˵P�L ��v���6��f�y���{�}	䀴���@�щY���:`��j��y�R'!�K��H�H��򏋹y�B|�|B+ �{�J��V�P|Sn�`=��.76���:����d��.m/��4����_�'_��a����q*^�-�@�l:oY�Bd�}�e�$�E[�ݷ�L�/ߠ|�R-�8ދ��?*��9󸂗s*u�ʿ�X���f����Ur�lʨW�mJ�������$=3Ezq-UT����%�*�B�_s��zt��DZP X�Ց(�'#x%��� x���"?����Q�\�b����VVe�v�~��ĥ~�]��qC���X������$�nG�M���V��ȧC�ضc��#���l;���N�"��ꇷ���n�G���r5�]�0���mCb���+"e���.M"n��ɧ�����!jlr�i8�i�����0��%[����u�RQ��<���%�1��ˣt��M�?S�Ʀ�9���h�E���0��L"L��3�u5>5I�m7.c�:"SJ~��?+dKr�'Y+��I4���:u^ʦ1��Պ�Ҍ��=h�\ʺ�i�B~�t}���ߧ����-Q�S$�=4b�O!����V~���&���?@Zԓ����գe���.M������H�8��e��� s���A+)QJ�r�!>��E4�C}3'��ը���$M����=C�7��0i���\'�,�+C�}s '����^J� �?�Dg)`sFE ���o��B�x�%$���z�����3tQ�Q�v������ye�X��A<�-�=����/��=l:6��|�PG�I@�1�}'晨wWѫ������R|أ�>�FR�geiՅI�Á3���l;I�å\Dz���PX(!�^ܨ)�/T��!�����&��x6Ֆ�����Yx)�}�'b��~4B������� ��XTR�Q0��Zξ�Xx��il&C/^��g9]�c���|�9��~�������N�¹xg���`l�塢�	�vN��LU�d��decM���r�I���k��Y�Wp@p�di�ǝ][k0�3� �df]��v�z�'408��?�U��Ĕ�	/�6���D�������dy�N�`�L���%o@{��h�z��N�����1S�@�:����g:���2��0ǯ�^R�s!_�ɒ�a_�4�9\��%w8n��<�m�U���5�d6oz�����0�Qh<n���������![���B�M���b�g&��x��ەe�65z� �4�m�Oǉ�	 -ܙ^�w��v�WkzUg6���/N[�NUn�<	���`_=%Վ�(sV���_��e�g�7�ɹ�J? aW5�*�Y�W1���*��J�C�sW-J�E|"d�4�M��ghG'('��s�n�ɽ�����:b�Ȉ�ޜrS���Vp
0���]fK6p�겘��Ц������z�)���������з%�^|���qb���b� ��XlxVHYEB    ab24    1af0/L��-��JǼ �f�S�ݺ�£A �#���[�v*�5U�E|F��L�ï�tL��d�;6h�	l�<��i���01�EU�ܑZ���~�0��*E��k�-�F4G<4c�O���?�H��rno�� aJX����$�5B|9�&-��aenx�0�m�KZY�9�Ё��=6�,�B��37��Lwb<}����h.N�����Abh	��w!9_nR����\A?"�v9>t�l"���r��.�ef5<�cPQh�FD;S[���v}�p)�O�X�!RP�ކ����9g�2�R�Bn���Cz�տq���^#]+))��fU@�e��ke(��am�wS��5�a��E��O�Q��])�1�Q�o�l��ǩI�I@mL��ַ�9��<t>B�p� ��"�f��ڮ��q*��]q��PH�����CK����f/!5���!���)�9b
��8���a�Ō�oɘ&�f���$�{����xp�Y�2�ɐA*|�2���f{T�_����B�w��I�p�u���7��|�tkB��h2�N�w��E�w����Q���ʟ@/ �(Qѷm���m���/7�@Ynf4Y�QlM`~L�ٮb��ln?�����|�z�N����~6��I�8S:�O�[��B��	!n�����Gdɹ/Zo��G���Č���d2
��V��X�Y�:V��,����F�K��Λ�U}�[���u�4�QJ�-��g�n�·�Ǭث,>4^h�P@Rz�,�T�wwX��VE��"�����(�dXK��]�p�5�Fb�sn�3�{�@g�X?��Vi0�D�h�[Ybf�Z�4���O�BPȗJ�nZnp�R��x��Hw� �£�\��U�j[��q����ha@sl�!+` �������ӥ�DD�Ii3�2U�Ǿ,���۠m���Yoɭ�E�y
F_q�����?�x�9R蛤ax(���
W�z֬��!c_�����@�7���Tڍ�=?�}ԡo"�x@kC�e��R�F�+�R�����\�Vd�х���A��X�r6���P��7B����J1u=�G?Kj!Z	�`Vt��R"��'��<��8_��=�Bz�s��$s��R=K�nK��Rf�DU紐B6ر��c#I+�4�B�n
TS����c�2�-����i�7�Q�Ͱb6d�@(�Pj{T��TY6�E�hϒp>+u�b
z�Y9����X�p[�l�.��z�͊ݘ�� V�{�5�*��'co�z[��0/�6Ф���'�ICGk��%�Sl{����28�?�=�*�g~bk�X���XX��fM>���g���t�@����v/]���n�6�`�,26H�VKrR�P�_Ȕ,��A� A�_�ۉͧk]e�yXRY>�.E:�W���������P����*�8�W��h�_���M5b�Zz���ʸYO}H3�1�E�ҷӠ�C��n�?t��"�|,��ڨ~�5����E�\c)��f��fDƶX��Sa��˓r]/f�$ر��g�{R6�T�/
�M��N��P֑ct7�I��Do��A*y�����곎7���"O�L�"� 4��m�E0���j��zV��[�4T��Dd��5)Zk���Z@fD=�R����V��]7O@~�U� �������`ˑ�r	��7��=�_�b-v�W����zz�����<�i��X5G��:WO�ay��bj�3Y~��v��
�6@4�vi�-:���ҿ��|+���ri���,�쐣��Kpp�+�U�@c�(�+j����{�W�%!���լqʭ�\�xWB���{��amѾ�I.Q�%W|I��h֗*����ZT9����4
�{�CZ��u�}�@ul��`�B���1���ܰ>�߾�{<@c9�W�逳��'�'/Pj���?�z��8�{�F��3�I7>�zk7HJO%���0�"�������e��0��,+�����zG��L��X�J����Q+��_�R�IRՍ���"��D��
�_@���s��򴁵�y��o�eP���|�J�U�6�v@���6J�3Ҷ4\�����[FŅh���BP@D-���F�_���:CQx0���B#B�R��`�;L��gu��{�n���
R��������ǥ��A�7�y��rOl��"��jE�Ǌ�8;є������Ą[+�kQ�Y#�����e��G���}�E1;U��-�.?-ی�s��@t����c��F`wm���;��eدJ��l"��2��=��&O3���/�A��o�������'eY��8�y���S�bm����b �_$ܩ8UMYH��� z�;��1�	�?`���v��ik���������/x�r��<"�S[p�,�ɝqRׅ�sqZ�rsl�IZ.ԲC_Xn/<���_%څ�a�qd��HӼK�}�wC�)���SY1��%��<z}�KM�Q�
����(.R
}
Ԗpi(#?_��5؛#�M�7�bOv`�7���W��x!�2WyS�L�l��%�+�j�n�z��9�э��>�ʀ��vbuP�-{JD=�Ome�#�I��ܑ�$E��dbvZ��*%ũ9�@�wg�j$|~��Zu�ʴ�y�(ِ����>s�p̠�I�:�a$�̽'&��(��Ax��"��u�I�?�iyCvIU#�Hp{fvZ�Z��M�G�AQ�����/�_d��i�QI����u��i����r�{̰�B&^B�eM��A4�-�7��3���ʵ������g�YI����o��`��`��2��{�_P�<�u�d�D�]�3���u� iT4RkGrS7���(2��z���.�dw#�_j˔'�Ց�h87��8��pF禛��[����* �^�:A��
�� ���H�l+�i��">�/���]�8YF�d8�ؘ<�GAqі�0sX>�L���It��>ǭ�}�$e����D.�1DJ�]l��۫f��#'/�Z����fy2]���p�)�C�Nu>u\�,�./�q�Ɣ����
nNWR5�ML�B�����dQl�+�ZSKx�kcΗi��\F��Ud$A�΂�QSh��Jc1�=������)�[�\�cv�W_�j���`���*ϸMD���������͎�ٝ@�K�6_�`���@�P�����,�ߒ�VúX����8��e����j����d��ۥe���U���:F6�c������G��٪b���
/�f���n��ba�fC��q�Н�c�s��9�v�Ɲ�)�� �sG]�#ly�x����U�ˋ�ɔ4��;.b��Qx�*�1�?]u�l����j��(i������/tX$V����"*�$tx�w�dk<��	��kFV�M�~�Y<0�<���ĺ;q����79��B�_�P�ze�篛�a��2�6�8�FB�H\�;���Y����c���K��Si�TQ�,�l1dD�~�<���A� ��Ryv�@��ս�a�����ZXo=u!H�D�ϕ�%�L�7���uT�<jF��vM���"GG��S�)�6����2�Ҹ]ݷ{����H�r~Q�%E�9|��Y6rdXe"���H�#���v~F\1�r�t��1��#K.P=���6ʿ��f&������9|��kwBYe*�I�^�z蚳�aPȀV�y�WB���2^��=1���mӥ�W�H����U�4��AO�k2a�X;��ا-�WM�$<m�l�Π^.��C���|�m�u5��ԁSkpeR�E���V�6�br�U�m��׍}�C�/�kv���g�-t��(o
7TV_�&���q�ځ,r��S�x`V�d`�!�_m��E�)�kMb%�^_�8�bz��/��I<�>bU�;L��ӎE���-=d��>8���C��z�����d���da��N^RC1J}D����4����?jHZ :la5�5��TAfk��i-�>�V�{��?� 0���&�T]�-��@]|n������Fۙ�1�R7�Yw�P50E��rp�9�j��O�c���G�@���e���Ҥ����M�oTO���JGh���$��f�$E�^��>�!��(���K.��c�.=R���o�p�|�Ҽ.j��J����<���xC�z�l��^b��]�wO���t�����4���6c^��'L��~�X-	��S�/tz��!��ol* ��5,Ĝ�B		�b,�ahxx�	}F���Ho�1�q�sێ��ýGj�2PgJ�?f�[�P��!\B����~3+��"(n�!�
r��3e��/9?����X�4�<|��K�!�ƴث�f�L>�V��_ Iq�I�	�q �^�8����t��ll���Y�Ă���ex�#h[K���u���s�*�M 2�B��e�к��#?��6}�Y�xr:֡2N�[�ᢪ�h��{W��_7�g=k;��S|��f�Yx���$N;�M��q��ؾ=��m�"ӓ��5�;j8U�x[ޢ:{�ˌ/�^O� ?�	��NX8ڈ�ӻ�B�ە୕���Z�E��X��c{�h���e�KS�,C��;�E=�br ��Y���m6ޖ"�1��Q�'�К�k�ß�?��ޭA��2B��/�H�m_5ihS�ڣB��h�ڊ���:e�]Y��.|�+���m��q�&����Tjz��oPC���Q�uL'^��`���o������tݍ��2�C-F��:�A�Ӄ-�x���6��!s�N�t����>Ԑ;H{[��~(�Ċ����"G��8&��Rp,��ģ�Ս���5�w��������o�_��.=��6�Nf�B
{��j�L���^xe:~H�^�Pc��Ѱ3�תb�V~�+yi\6���7A�#`���(6����C����~<�\_Iɳ�d�ڜ�t��j��u��c[�S�_�@	�Wk����*�{3߷�|T��ρ���X�#��S�,[^DMk?n�M���D՛:�	�`�|��9߱����͖m,������w�F!��5�G�h��������6�GMd�`XWs��`�B��Ҷ����	EO��t�y�]1�e�0�H��.ҿ��D��yex>C��S }�?r �F *i�,/��E���:74���	7SBG�҄�p�Ű�&vc���(>/���0K����������ׄ��G�mG�����IO�X���iY���K� �#��hƷ�����`?(䣏T�	Zw�w�o3rٽet]v�Ԑ�W%Qa�R��e'�h1�4�u&!9�,72q��:���>��@��O?)�����b��j�u4"�ߥt̻`Nr�"r �e|��.�k�qRk=3i�	g��Ӛy�`�V�7Y����t�T�"����t�~T~�>���7Ȇ�h�N7P���Æt��_td�˴��2XY�k����6���?ɍ��ko�cL�O�,� xRj��rI���q\�f�)������B%(�.^�Z�1���_��XD�X]�"�D0��2.]k��w0	#c�JĞ��@7�E9]L7��H�����ѡ��4���b�f�N6y����3�+UK�2�}�,?��'�^�R�4��
�ρ���:Ft���oV��_P���
��ZM��	��� ��N�x�����&_Q&.���u�r&���P*3�YrZ�ŭ�>��Q�Iy�n(w�$>w*ْC���Z��|Hs��!yM����gznܿ�X)`N5�nM��\x/��+�JQ_�k��x,�5�B�+�8Sx6���i�
lB:� m�-�-��������x�9�8-��ܿv��вߨL[�K�����IU����� ���vל�%�)9(ZGj�gW5�ץI���9��Į�:gn��Ct�|��>�%�x��)�ײ��B�ɖ�gyNt�I�z��,Z��*w��y�\%�ԫsz�dѰ�� *6{ioЭw�|Q�_:�;���TG���3�6����h��T����O �����1�ڲ�g�\M����`=�ŉφ~V��Qɧ���@�f�}��V�����n6�3�QМ�#8�.!���U)¼��tّ�5P:����!2ӹ�1/���&+o��ݕ����D�)�]�!���wVz�6��Ǣ��'\P���{U^-�P�ɋI$A�
��aoU�5)�1�5g�EF�k2�گ�B\���|�Ѿ�o -s/�`J4a]� ���^}B��B�fLtI�$g5��x�yDeuUS�8���8E�Li�W��UfHF���'��т�����A��#�p��dKx_��Ε�=:\�c��;"x���f�#F�ٟ�� �$!y�5_#+�{io~qB�\-�F��3���7Z��K0PƸD'�a�f�����u�]����R��wº�M5����0��,�A�T�J�Ol`D	��T gO׀�|�q�Qfր;ʞ���g4CQ����D1���bԊ��Bv�>[�`�:�ߴ�P�*re�{�7X3��@c��e����b�H0��W>:\ߪ��bZ�����m����Ӗ������i�_@�89���O�5��xzD�/��Q��B���Z;�5�P��A��TpU=��!�R�[��
�[:V�E����2�i�J;��	�qξݜ�*PR2zn>�#���xH�jD���N���= �)/�\Ƴ
Vo/@lq�GO�i�x�xK_c�Z������_�=����v�N m2��b���ph紀9LO^��â�.5�/�䞁P�R�����Q9u�X��T��V�JO�+	7��!ۀ3����(�v,P�Z����f����Q3�"��$%��@Q?�-��i����_�P�����e�'7����^�	R��c�N�Bq���˟;j��V3SG�k)
XlxV65EB    2aa2     b60GP�{�~-z����#��"4�iA�Ә(,�U��Ply���|���5d�U����k>����3�!�'9��V�߂\r����fa���86@��N�p�����a��	�WF����wp�[�6g��nHьY���2>M����1�kOJ'F�Oe�n��QS/�S7I.�� &28&u��c������ 91g�ʭ��B�v߄J@%"f�����~���pc|��,�E�Ĺ�OC�ƶJĝ���) �i���;��:8��/���U�m��ű��~���TS����z��QQ2h���!Y��5�L~�ysc��>rd�y�0K^(?H
��`��{��(p�ʕ�= &�^���L��i��%\�eYKuQ���u��xΜ]$R��y:v�������!sa4��+�cw��\.ިB������y0�R�V�r��6�p�����c�q�9J�aAL��`�'��NXb�
�-��0F�h�Z�YY��O�,��/���3B�ھ��?��r������掗����)�`R5�]��BZ4K#c�ώ�e�C���F.�֞�y� ����oubg;I�f�����=�v��Jy��=]5�F�V>��A�E*Vs��1�#8�3oΊS�'�ZB;a-S<�!�My��jS�Xv���j����wf���3 6J�;�I XgUx@Nó*�E��B�����G�hg:m;
�L�V��_i|�;v%���2𻬵���6Oz�k�����W�MI���ޯ*/b?�Mj�Pҋ!��N@��seg��d���7��{4�/�k�9�d����*6�+Qqv&�� ��.�#;�괭I/����Mzu��Qb�ߍp*�-R�]��6�,qR��#�Y7SY�z����p�������I�D�RD�C<M	�`k9Y�.�9��+����d�kɆ�dɽ�b�AW�nҷq������̴^c��$j�a�/�L���]k��G���c���� �+ ��WJ�I^�M�'�m�~�㞜}��x'�p��\qk��"%{,�9�����mvr�U� �UW� ����q�hf_	S5�IZ^&�W�\6�ϼ�YjR��F���l����.X����91[�aਂ������U������v�����%�D��%�+ǹ�ǎ\O���蜭�ڝ١$$���dJxQ+����E��P���Yq\�EO(|��|�lB���J�z��w'�!>��ld(��%���6��<�k�g�֗�|����'��$dI���z���˗���9����i���\��W3j{:N��v��ʰ@<-C�����忛q��}ԑ��
�L#O���ap,���ezda��(�$#(H&%����(3]|k�6�kC��E"�]�v���l��/_�dW�c�$��ݫ�z�,�@�JuPie�2k`��Y��<���{�_���u�$������E���`�]#�������񃄓�j~���J�R�+A�Ԫ�9Qǣ s���{7#[L<C��o�R|OB4Բҹ<mu}Nz��&v
)�邢�/;���p,L�Me�٬�3�k	"���H�n���P?wߧ�Ros����*:�!F�Є��Q�|Jhw+r�P!]ߕc��6���C�P%��'���\9q��V�G����8@��K{���KE�w���B&eA#�ȜY�kU��EUw��Y#3�(*�l_�,Y`��ҍ:�Dy$<��ṃ՛D�y ���o?��n�����M�IG��w̞�l/�+o�6����/��u��8uH�	c I��EM�T�h��_[u�o��y�?27������=���E��Uw�e2��ʽ�;tT?�jn�bb�<����0��Ma��{X�h�ǰ�/����/>�LV��	 ^[-��RۺV���I�4��o��}��.�ҩQa8�h�w����6D���fܒ��X����*q[K,����29�,%O�A=�@V�<AI�Wz���[fւn�O$F���ց��$��ٞEdi�2�q��n*!
*�1xԧ�f�ń_v�*�,��E�*�&��<
j,+�@W;���˛�9|I�Pv	��J;� ,WH�r��=Z��S�ը!��I�2�'��sM�㎚���C���e�jڼ�(D�֦���	� ��بrҢ=gh�!`?���'�P��]i���3��a���L�'���r��h���,��E�0ݹ'�:MI�Q|�
��n��Gu�F��]_�m�D�F���H���y�)F��
!gx/�X-9[q=9��i��ݪ�뤒.�'���0�|�W}�6�S����/�T;Ң}�rO��*BE�K]u��Lݍ���	[�I
!�Ak5���<H�[��R�@EO��̙�Ԏ�;DՎSe�=�g�#��D�����h���_���L&�`�P�����,�L��{DQ���պB�P؛���~K:�r5d��b��(�X[Z����&�B%Pi��wL~Y�����Mzo�����t��^��}�t>�~�,��rP��^�}	�E�����iңrг���+�*�`s/k��R�A�q�u��8�/��Q�����,���ᛣ�Nh����C'>�ى��y(RS �9�cv
o�" gba�UE�oK@4���^�'�Y�!	�l�>3/�42{���e�:p�+�.��4�>�	>'�_m��Å�E'��^�J�����i�7�v��d��~��OI�E�#�g}��A�k/ln��B�y�ћ�u1�4�V�T*�����?'���n2�ʏ�O�l��)��z���%}�Hѽ���B�.ߗ���;:�A{X~ߐ�\Q���.��'ۥ�b����B��y�<y>����� ��dܾ��G#T�h���^p��@��J�������8Rp)�������a��s�8�
XlxV65EB    fa00    2ee0��y�<Fr��bƴ�dMx^�.p��GףRjv�9�B�(����>�{��Ԏ�C��{Ub��p��j���s�H3(>{���a$HVU;�����E�$aH��	Ð�WE��83�?��&m��ޚ�ɚJd�̤��J�uNt�* ��۸��W���1���(���,��<�t�����vM����3 �kc��������ؿ ����z(0 *�����S������J�X��t�EZ#C)������˘�a�C�����7l�w������ɓ�F�ޗ�;9�%��6�Tiy�p��1��7�RJ:B��gt*~��]��5mbX�nD�[[� Eu�h�M5	}->b>�j���G�w�w��ǻw
�ۃNe��80�i6Θ��/#d$� $�sbz����<>�������l??KN�+)iB\ʙ?eL�&��
�*�$d�9��!�d�Y0����1���C�~7��Z�0ġ��H�κAl�z���WCƋ���+� �ֿ��۷�2��Ӵ��fk�����v����|B֫q��ܴq�	-ƦQ	ev�X=�yv�����XX_ݮ{��B: ��h�������E�j��v1]CZq��N�c��|����Z��D�+�o=U�\Hl�B���u�vo;K]c{b��q��������
�/��J� aK��:]F�;~�ࣻs�9���!2��Y�2��4-�S.���CS�HY��6Oo\����%�Ia#�L�$��̡���}�h/9�G�}+Jw��v�m+�<C���f��{��\�m�T���v#�����T�U9a�=�_��R�~���	.3y�ՈI6�B�f9�L凒U�n=H�vy��P7+��j�cM��΁-ֹ��)�}c�s�Gc���h1���p |�@cШ[�CdS�MB���	_��CN���"]�콧�?,�[��EX�{4|��=-ہ������%���^o�53~� (gl�VJ��$���� ����ٱc����k(���/iF,,Y��苶�YbʥN��۫kÉʡFMc��K����/6���,"�yC�U���º���6��q�D����5:���4�����S|�4�WN�M���yHD�pɤRZ)nj{Ֆ�`���}4�Y��F<����ݽa\�g��%W�J�:�L��є���y6/s�I��q� �����;��TB@�(�R�,��,>��PX����!��ɘ��o;<M��y6�O	i��R���L����k��)�
];6�G ̊�i{����=4F��,�)�i���>�&��ӓ�l/�T�����'BK�p�
b�+�{�N �Gim���7�8�'�lsH[�}::Qq���nڌ���s[#0�e�@4��[�3�E���K�WLY�v�	l�����M#|}������@Ÿp`��uf�uZ�H��\d[����_��Ը�s*�0J�~��O~Ab?ɒ�-Ԩ���,�	��A�A �A���L�2�De	��n�}�^�ڲ7W0T��_���cY�� =�r�=z����
m�iD�I? �&K`o ������i�[s�ʾv�¨���=����S�d��@⭦���uڽ#����Ƴ�X)b��21/�B	Ϫ�:��H�o_ZB�!�rK|p���)e�0�+K��{�>ߌ�5�8||�wC�xX�rj>�4s�a"�G�$',�Ǆ��T�eT��'�s*��8T�a�0��eH�/<�
x@n�I� ��l
 �
)���[I������~�3�,j4T�A\s�Z莶<�P�6u��q��h�f9~�;	8�� �+�{q�g��p;7BG&s���ݲ�W�ת�ILky�'2fU�P|�.�9`j_�4���p�']��6��f^m�P�qÖ���n��1�f����]��7��m���6u�2z�/�$�*H&���䖣���I#�����q�����������.�ɯU����o� ��w/�j���q<?�Z]�V�]��<\�sbj��Ux�DgG���%�#-Z2��(�?-��:��~�L�������c���0F49�v$^������\@h4hrОҢ���Z��>��*x*T�"=��0�ŊUK[���ļ#���{@�\�|]���D��ZO���s����kkY�g*�:�h��i�`�����-JL�] ��t"u$�+�'b���zJ4�AE�Uˎ��7�!+���!�3=��k����9��ǎ�-���_^�\��l��v��mb�wp@�z��p�
��:_6�}��nR˼�bE׻C֤3@�$7<נ:0Ѳ�vE9_8Ѳ�4�k���ђE�<���||�Ѕ²q۫>�<'���p=2��gH_��P-\����Ņ{�����L�cf)x��&jQx�����Z��>���|�w����o��*J��i�����u.��{>^1ҁ#/�1��>%)䙘�d���M9�)��f����.������HR�ms�>�)^O%�Sg�Sm�H�L�cR���!�Ϩ��HV��z*�g�(��Z`ԉ��iF��np.Z	ޯO��"��A�6"�4F�Q-a���D�G���3���5�:�@E���߃��j����t7n*�����L���D��jEZ�����p���&!���s7Ɲ=�Wë
p�cG�3)�g�J�x��Q�@  �Q��J�G�v�9Q�&/ ��$Hbۈ����Ԩ�!��Z!d�[�ܓ���
��^a�ѕ:��e��ǭ_�q��S�W̽��wĲ��C'O�c�At%с���t��,K��z�V���	+*�ϕH4��"m)q��*ف�Z� �y�B�R�~�M�㸄u{͓���7���J/zQ]~C��9=��73Y�IX������t�U�'tW����*$]\
h� ��$�z����c�˅�,.G��"����~XM�lXB�.�4�G��#"�c/�혘����Otm�y����5c������*}),�����G�+��"X���@x�����P3���o?؞
�7�@o9��\��r����WF}]����:cf3s���^Ȣ��Yz�SҚca:w�9w��Gt�s�
ŏ!�:,ȝ� .�es=m�B�\��?����������9�C�} ��F����j��D��5�@�~Soλ�6�`�V��H���Ͷc���d�x�`Ư���ʛ��bx�:fMF8+���>Fݯ�g���7�v�k�;����v��T)��������Ð�[� T�A�V�|��o�Y�3jkl)��B��3��B��*��y2=lR:�!d f(?*l��+QR���Mx M�D&4�6��׌��rC�L��PyCj���W��s�»-f8�=��
���3�&�-a� �C!@�����(2�o5I���ý>���Gv��8n��K�)��hz;�2q����0 ��?3z���t4�Jڭ�7�4:� k�ʁ�3ӫ�[�[vԀb�߄���lE��-�t ��iqf����>2﫠uM3�&D^�����ʔ�9�G";�F�iq���i*y2�Ĝ8�6p.������EO�|���i�q�>[hO��&�꤂��i�i&m@�Ⱥ�N���Z�x�S�E
ωVMQ<5&G�:Rs%�Rs(�e���(���D��w��0�'N?�oR&f��V���/�\1<�;�%e��]T>2���[ac���h�gK��b�z_�}�H�~Cu|�n���9t�fm���!�:�ϏaL��q.a�ƞ#���K&�<_�R*.�t*�8�V���
 ���0V�չ���Ԉ��| u�8n�q�Fs���V��f��*�GM�
��<�s�&X��-6����֣D-��.��2�w3�	�������|u�"|�.�����6�&!��	���h�������nl�u9#x�>���G�$��N���"�Cq�e�lG��3����Z�G�V\��'��DB(��-_U� d������X%Į@'q�U�ۈ����\P j���ܽ�9��mR>N�c��Q�b��;C�vqQ�M!I���ǌ��g����y�eΑ�'`9i�_��Et.̄[�*���*PA_�{�'����DW����3`��g�IK8rp0��0�2�5�P�Y�E�^��I���������gJz�	��݋��eie�Y8J�^#C��\pJ�>?#e���:��5�dIr�2�a��b�ȅ�o�ӧ�`O
v=&T���2^F�5OA��S'̊��u�5�Wy�\�q�y[rV��7�Ȯ}�b�^��o}��Y��X�@� �Ǹ��΁�U�枿��O��A���H��Q=�m����^�7�W�m"Z���'W0i^���wg&#��~,g�"F5R,}���وyr���]澲L7�i���^>{��,i��z
��")�jO���\��ʢ�<�������A9?�k'��5�ǀ�w��Q���"Rm^M!vc�'>ڙ���wQ�wLj9�_�=�_��
���ޮ�a�C�����T�q��4�"�J����j�w�Н|E.�I+P�!r!��)ϵ(�G��kD��������B迤� �Yw�dע��Q�����#c��������;.����sc���4�W��P�ܡ��创�� aI�>������zEE@j�V)����D����� �{R��]�=2�����9/�̤���} �C��e�6{���	�ña��t[=�I���?��X�Ͱ�MJ?�����l\I��Unc�#<��R7�mz�ެ����)w<�Ϥk���Vt��i�6ү�����v@	*_�$1T��=��
�"S���@�AJ6"ht_q��{>��P���籋����#�T%=�P��$�O?��"�%V�o����'ULCk�����<�Q�v�K}�m��/��D�0-�vc̏./M���L@+B�	�C�ւN�!8<�`�oZ��m����m�?�=Po�� �p�r�AE<vS�8`�\�vD������ i���uߥ�t��!�l�����f3F�N�B0����6��	C�U1Xs�FB+%t%1=�[�[��S���֝#5V�_��F�����uL��G���lh�Wb�3+�/|�."��������)���\L�2J�i�����#�q8
~^Pzu�au�n��R	���Õ�G������5>���QJ�I s���`�u�6_����[���S�F�ߚ��Ŵ���;�Jj��i�o9�Wq.b�|�L������� i��t��c����EX�ٞ���u)���7�F���q_����5ڡ�0IQoU��O����k(�8���Q1��p#� H�A�`d'�� ����aK2�v�Q55�?�N���B�y)X�9�np�3OM���품kw���3��)�ܻ��mPL�^g�N!���K^�,��=;;���.�{f��	�����,�eu�$��u��5�Aqe_f�>����bz�|�o��`�8d��$e}۫T?�t��u�Ov�����	G=m��f�Uؔy�զ͵P)}&���\����b���G��)TR����P�C1_�_S�0>SǞ5@�b|�a�+��y�`F�T2l��� *�;���r%ʶ,�����L�[F������E�Z"d�>�Z6O֡؟��`0��M'�J[y�PPQ����P:���q�O�^��~�~�;ǎJ����4e�L�6�faE��\¼�f�$tt���8ozHr�;Q�N�$ߩ4��-����`���������lzpJ�ZlYo���\y���h�do���}c�B���]�qF���~�R�ß��p�D��y�&O\�vUg�1�Ef�d��_1M��t��@$|PDv���M���^�����ؖ����_�4B/��H��3Ђ��<`�ң:UU����+!UVD��D���%`W1��AⰛ;�d �W�##�~l�8�e)�v�'Y$�̬+<?�鉜�b�Y{�4�O
<a����E4���p\h��wf�s �ɻ��X�K�d�L�K��r�Ƀ��}��.?]�hI���������0�;����|��	�K�l�H�&���4��F#��z'���F���H�`�v���W~�[(N�mA&.�e",܈]���R�k�B��ǧ����:��Г@���K����K��B�'�[ڹ�]=�C��Q�T�c��sw�����cV�E���P����b$���V��^5@��>QJ+��[^�v���>��~aq�He�l��U�[������s�`�b�t���πPx>�ir#�	-OK�p���bG��u�}��,�7�{�I���wdcJI��>$�N'
���W--��*a����������>��u�!��ml�|�<�
�h�n9�r�.OG�o���.c��w�k+H^g�p��-��u�p���h�F���_�����Rx��/���2�
7��d$r�(�N���N����|8�Ζ¬��(�Y鈺�x8<�f�H)�hx��v�L����t_����e}Yl��H���"��B�7�T���Ӓ�sw��9��8���9���)�Q��ZzN�c��O:ˇM��㮅�½; �e� �Q`���B�!��0���4Ahv��������8>]�����pr�s�����~�Yq�X5�y2T������-a��&I��V���8>Ig�ΦPx�t��e��?�������̙Y�~�n��e�V*W+��-�J�Z7�_���[\��Pܣ��`������' ��~l���˽����z+�yB$s�s�[i�صԄ���r~�G���	�7��ο���:�`�Y��e_q;��\.V���\��3�QT�k�v�L����
�G�Eœ���a�J<XL�k:<�2ـQ��dVw��g{ k�a��dM�Ȓ�6��?��O�Z���ᐋ;իL,�͵��_W^��9лr&쵶��U���VNYSn�7:$��_�|
o�6�~����Z�b^�J�s-�Ɏ�u*�Ul{��|ll������޹G�ȩd�Zk��x|��q�"ztr��~���,�ȹx{r��k �� AM�Y`���`G��_��_?�[Ew%8��%���	&�AI��*��*�}|�>����n%C���b�P� ����}�
Q���e��6����(�c���t��ZBk-gڇ��2io`ns�F��	�(o��ޮl3�fC;�C�K\L�ڎ�,�Q�.�̢P��`���o�7�u��'
��sbP>�<kً������i��A����U�I�4�=9&v]�5v��H�
��y���>��&*�WoB���@;iJ�����ֺn�r���E�i��'l�G��q:zAa�Շb�$��x�;k�>)�V��쟩���r��;�h xA����$dbq�����i��[��O�J��COF��V�c{�w|��{I����Z#F��T������0u_�H��3L~��I�;�ts�o�&t@���Z&�Km��]T��V�V1g]ua<�'ez��T���8���'�zr��ev�����]�x�&Q��G�{@��p���ˊK��jJw��zڡ�>�g��K�4?���!=Sv������2�=Wؗ�~�-X�g��e��^=Pu):���b�`=���-B�51�>�<�R�e�1G͐G��It��D��[:�i�䀷�V�C�NR��E�_��2����f>�/�N3@WCH�'���z��9�����ܐ�2h�h��O���A�>u"����"�t���|�Y�^�24�����:���^���Z<��/o�I�f�L��dy6�ޭXz��@4���B�Bm����YZ+���!�'��H�?<�*aJ�¯V{CC�a�?&q�Cd&H-��q�hH)sT�k��-�k���و&��oJ�#��sG�E��s"UMU����xe�E�qM!�}�h�v̲�0�N�4�e�g�j��(��j��&"��	�X9!��;".0X3
��W�_\m3+�����a���ņ��>Ў���z�䯏z�X&k>u���V�3�P�\�y�n�i�����'���Io�U`�8��T�ք�G�"/H`���R7��^��AN�!���8&���Yċ��2�9�H v)0|��<V�D�Y�?MO
Z��qA2#! �fH��;#������f�L
�Lvy]�0%�P������_3t�*�ߘ	-��=�'�,C}��ST����3u g�qp�r���&`
sc"��Gh}�1w��� �?�;)7���݇�$H*K��R�J���|N�Z����O���P�Oųg�S��1H��T��h��R��=��Xח��N����pdQV�p��Ϸ����=�Uk��a9"���	��K�����s� ���߄�G�,̙3�u*����l�Eh��?���-�D����ex2������,)T���AS|fx����'�4�����2�(�1p�3'��?��?D�!lz)�`Ɲ�{#��F79eї2'��n7x�T4ot���������&䗾�r�Ѥ��je�#r�ĝI�~�����B���#n�f���Rt�n�~�m��y~&�ۇ��?��7��A�����b���)ݡS~S
c�2�A�"�/�RI��qįx�R��jX�1�E0ڂO�ID��x d�VD���g�f�s�ѫ�K0���6}���BH��$���m��S�$I�(%�(��A�խ/~�[(u��c�J@���/)o\�E����q�A�-�S4�&�p/�p@�v��膀��<Y>���	\�}�LϢY��_��-�ND���S�����rŏ�逧d&B��I!�qnv�cnǫBԇ\��WM��d�Ps
y�H!Z��ҥG*3[|����Va�]�#��#�(ڙ	������슩e0��� ������T�>��M��=N6��]o?
y��.r�?*��Կ�w_�&�G�5�=�7H}֬��'[��&��p9ݓV�����K��'�*���м7s��}�)IW�o���嫈i-��ʻt�~�=L%��FE���������@  ���)�o0ҿ�QT��'���O�u9�d�S��kv�q�j����W����ծW��xn�,6��}�L�Z���-�  �<BjJܱ9�րX��m�JB3do�.�6��(�qF�yB!1�ƼlӛD�p�k��o�5T1!�[P��tBf�5��"�uL��\ط�_�Lj瓙�[՗�5���g��$�@BJH��Q����1�	ɵ����X����0jہ�"Gb�o�K�V�q���=7v��z,�y��ϟ�s�5�y�~[w�������v���LM����k���̒^��zlw W߯������$ ���X�쐄�[�	U��Y0����~\W:�a�ȳ�]}�f�]���lx|��Y�}<��0�Y�c��D���x����/���ȗ��R��`�<��'Rq/��c<��C��u=U�I�PgX������鰻�n7?�7�̰�ALoofh:���7!�Q����q���׶3��֏ƺ����O��U 6ʹ����c]��(�D}�8�a�.���FDC��\y�w�Dgw�!˥�!Y�+k�����0~nG�ݫ��d�N^���3"���\�@�M	+�vg(�``_���K���=T�@��l��]c�]��8?��BԢ)�h:Q]���Q��� �y�v��РjI�?��qY͑k��{i#_�d{���|�aX�%��S�.���}N����9o+N��j���nr����r��Jk
��xIX^t����|�,�YN*��i�Z�Z#�B(}��/�.09��wp�˖��,+q'��ev�F,]���0�/��)OO���6�Z�F������ʠ�~c6����I�[ �c(؉�#�����\Q��������T��6�au���]�]�~�x�L��lwIͥ��P�Na�L�ۋ�|3�/�`�;��I�
ކ@���1�L���&曍eU��o�����u���@?�S��"���+FUJgoM����U��(�����i�̓#\���;/ƅ���	�D�?��#%#�6�Ҟ�&I�A^�i���/]��1C�1L���hNm�[��[����_TP6�������c7�M�T������g�Z-������)�d�A��r|?b���~�:s��p8���KX�������`�S#:���t8��m�E}Auq�j�����!���߽T���=;��\��Qݷ�VT�}_ΕA�I
��6�i<3=�	��ţX��E=Ď}+��Hm����Q�8N�3���B-�&�:�A�(6��3��p�:���2�ɀ���	�UU+}Κ�
��Ԉ�^�n�Z��#пFsn>wY���6�{��bR��{��!���z��7P�zZOV�ڜrݖet�?V/4o5�r�Mp�'o�TϞ�9r���{�G����~�mE�DM�I��(��O�g'⺡d��Cb��*qJ.���b:�؋ga&*}S(�BQ=ۤn�
�:��e�=�C�����U�B��.�Jwu��O������`���;-�^nQ<ٺ氳��^��f�+E�9{�����"�;@�z�w��&�I$��;2oGWV����>�Q�!?���.;&��-������ߨ��f6ZF�(<(����c�\'�m�����OqF�]�b��.����Y�Fص�������Hbg	���l�d�׹�#{Z©�X����xk��T:�΄b�+��#���� �d�i��$r���)�h��C�tKz̦)l�a���±�E���������o�?��)�t�&;I<@�h/��E�V����Q�/�a|�(���M�5�k"�	�_��U%��x�_C����LH^��Db�T��M�F]�\)��9��3���� 3U��s�:+�։Z28�f�& �/��[*q���Wv\��PdU�]p���	�5�j�v�����;D�AQ,��꺽9z.���P0�����醃ٕ���ib�n��׺2�2�6�iyȱG���]�U�(�A�5:��ˌ{G�6m�K�m���P����s�Ԇ��B�]�]�l
:�_����Z����x��1���X��#EAy�M@}���:�s��ϗ���n�����
a|��u'5Oo�s��wN����#N6X�_�`G�ε �tG�/D��J��y��!�ފf1�u��&�UB�����--4ٲd=k[�t���+T3�5�y?iӢJF���N�v�W����D6�����\��5�r��䎐�@�j��%�Q�O����Yk,b������<������J-�J�Ɲ�v�߂+�6z���:������/���N���A?�="Si�J)U��2
�K��-����'o��#�`���tNn�]���V�7Z�l�ּoC��v����M�Pz�Y�  �E�@���[8�#��Z6,��0�(�KƁy*2،_�b��]�r���q��'�z�~�e��qQ�!P���iO��eǬ�Q�vEz�O}���ZݚҏMzA�%���=z�֊���fܖ�|q���zZ�+4e�y��*�"a��_����H�X�
ɰ��_t�Z1;�g�2����7k�5)�5Jhi�,�'���]�:re:z�IN�:E�M-�~iZH�%����JG��X�i���2�����q65P	zl����h_ZO~��J�ɘ��x㟃��W�O}�O�J)ngz�w�s�8�ɔM]��4ˠ��sǀ�L�P��Ɣ�p�W���wU�����?=�����|U]��zؘg��r�K��o�K�Wu�Lk/���Ū���XlxV65EB    d1bf    2170D���#�����)B��GF�J�����V8�JU���%n�M�t2�9�փ���hJ���eK�h�H2_���e{�6�cy=�t`��&����bF���O����Dc"�U���?�O��Ņ��~5���#��	�@��"�,U>zP����6���^�hYB���JO���ڜ�a��G�)B9�Um޲fQL���1�Ċ12�6��#Ƽ�zP ��Oȯk=�����*j�.�~�t�.�>�
f�j5����YD�FD���W6� <R��ﺓ�<��\�G����$N�KN\%�3������絗�BQ�;��T�S�-S�8\n��'���x��-�����f<t����ίeP�����3��0&�I�Va��1o;�%om0���2t���&�����b��Ӿ��t�5US�˺��� �Ĩ�¼꺺;�ˬ�f��Ʋ$�j���Ue�A�y��{��%�с�Iw�ȴ�|}8�h�vW����X�e>�m��!�3m���uƏ<-���$���l���fr���X1i"9k�&��O� �5X�˅� �&��0��ux���ה���0�L:�^�K���`���9�	k�L���D��}�#������]�G<U�+��ٔ^[����Grw����2�Q��5z��5�#Ѵ����H:B{إ_~��@�}9����R�+C"7I���Ň�/�kun�*4Ǫ�M���jFz`N�ŏK��`o�-dP��B�^�e�T�WK�[��9_56������P�ch"&�;�O� U�<��RD���EL!�kG��K�����-�5�b;A�"�ӳ��'��l�z��[+x����S��s��Q�U�[����8���J1c4)=����D.]�\ל|�g	�5�O���H�����^���p�U��c8��U/�9�Jh�.ֺ�5F�a���1����p�EZz!:Y7�Wg�h��<�@�a|�c4�T���+�ɍ�whG}��+kK/_Yr��V-�FA$�O������=dƶ�'0�$�y���~����W�ٜ?l���e��H�tM�{u5�
�����z�%p����^��vď�ݰ@$W�d��$��P-x�6���k]-1$�Xoli�������[<�?Nw�&�TV��H��7�L���ျ�s)^�u�����^H����s��w�K���r�W����H$C��I5����u8|6�χA��{�{��X�u��d��}E˟�3=]A�xc�X�2�T̔����IS�a�=�&7ӑ�+.���W�ܣJ��e���1��VT)!��_2s�E�c�.����'\P�jZ�U���Wp%� D
�3
uF
	�#稅0H���@ 	A��Lv�b�RS�T���K�����J�Q��r��|'��m�wr
��׹լ�)�7Mn+z�qj��K`_w\24ׂ�K̲x�k��f&��Ȫcm�t<L�L$uAI]��e[!�I��}�Wk�h�S�_�g�7�Λ��%y�Ǹ���I�(���(��s�
B&P1^���B�4B��:q���z��Qq?�K&R�6q{՜���r��c�#�J�A�ڪP�R��!@��]{�}��􇶔�.+Wm��a�>���������k�zJ+�	oSyz�8�z��pp��O��e2�����:&	]-�<"��B s\y��3c�����zU0TD�kA \���;�8b�R��_)S%��ё���!I�
��; :����F:����.��,z�yt�]��g*�X#�B�Z�%Y��x�9$�6�ڬ
�M4�^�;Af�s��M����U⮊��(��2AK���p���'l�\R�Wy[Y������#\����� ��P�L��4��Kʹ)�ȴ锚j�����8��cѠ�@{�9�K�&f�l�e�>x{:��`�8���%�n<��Zl�Ĺ����3�Iz/�A{禶�|4��vx3/ �Τ���C%.�&�(�s�c��дqʃo���X��J@m�Fe�Qo�ۗ� �7,c�+�5�S�	��ݮ�X�<nYS�M��A��g��h~<.�5�?��'5b?xĉ��h"c0���J$��_��R�s��5�݃�����ϑ��zϡvLz���s�ú`��:�/-��}�Co���8̉�^%Ѥ��1�D6J�{���'��#��8H>Mą�<��P2���ƽ��������(�L7�u'���#􏯨���yf�E���(4�r�>�����5m���\�ea���'V�����Su�1��?�e+m׻	���{��.>��sG�VQ�êx�}NfB��"ǟ��� X�ZԳ/}U,d�m#���q48�Gc淔�*�-J�\D/p���0F:v��*�����kyx�ff��a� �9!��s�,B��VO����3������.�JH:ҏ{$�t����d=�,�p�:Q���_�Zv�CD�������NűFs��:~��o��Ɵ��^uԍ����"��ﬅ�}�u�+����T���AN%i�~�S��j���'��6�&H]X�J�����6;Ԍ+������1��� Q������:@�w���`�v�V���@h˦��!NG-�O��b��n���q��
u��.��������c�Ϳt�j�%��했�D?i�+�PHY�׌��!��rv�3�r6H{��u�&�}�1s�6�:%�~~�o+��G�����v��9v)«��i^r��D�RUv\���E~��w�̆GQ#ae�Sa���H�|�Q�:I]@o)�B����%����>�oXK�ʂ��P	v����h�� j�4���-]!	i�-�1�oB�l7'4'U<f@ݜ{�>UhR!�6��6�H6OR8{_zi�g�t�ѶP]�p0��f �P8��{�)&��&=��{�"R��/C@Ֆ�Kk��N����qnچ,P�}9bƮ j$;�/�uԘ.��)��csp�6���=����w`A��I���A�'!֋�G)Zd]�eBֹ=Y"~���������;�e�9X���R����_��U6��MJ�?ʄ�vԱv��oh��x�-���ٴ>���|�vTֲ�����W�� `3?:�yؓ�	G"'���?y󢑯���kI�c�F
Z����^�V}�-^1q�ʫ��^����D��E�@���\F�T���Zmz6���|kr�T]"�)ݗ�����ρ��l@�b���8��I�ć� ����N�u�6����w#���Q���
Ո��eelh;s����|�5����6�ƀ�*�,T3IN�x)_Q��s=��tA�=
�0�¤�;���$��M�MQ_�A)7��f��C�O�2(%�F�)�����r������m�y2�PȔd�f��;m�~{��1�>�}�N�����#Q��s �p9�[t3A��ij$��`�&�j��5a��z��ۨ��.�wo3�T���B%T�`5T��-F��
���޽'���ً�0֠��f�1�OЮI2���2��`��M,c���1!�^UY-�L���E4�N?O��W���,�U=mʯ���w���Q�L[�QrC�b������h>r���{v� 9�I!�70}���Qe��@����L�嶝�gc-����sѕp�.�3�A�7�����N����
y���!_/�K�L�WǑ�!�^ S80���a{ OM�5 ��M#�si����
����}��cd'^�WᘥS�Oa'P�6�3f���<g$�͍Ԋ��d�;�b��$��d���wQQj^T�R�h�ӷ>98S���w�Ӣ2r�w�X�^ޫv�a	4B�f��ֻ=d�6`��e9L�sA�f�b��*���|rm�Wa�2��N%faR痷O)G�)������BY47�w)��W�x�>���t�_c&1��F�$*r�(�G�j}�z�������<����-ɶ�󋧗6���)����6�<�Q�)SE��1�$l�ܺ8V�pJ��i�ĳ�{���1�G�9���w&*(��,���j�^�L�݄��/���#m�˘�<�e`2^f��ڬ��۵�Y�8�Ѩi4t����Pǧ�9;���V�B��Ә,� Y04��M^�Jӂŕ��b�z4;���Z�ZM�����IY=�*z� `k�6n������j��w|����i�D>�R�64��!�HC̯ho/�c�t]D��z 9P�	O�{/A��Rx��"痪��j�rhmjLD���.j�����e��YVr�����pm�T�|J�8t9։����f\J~��;���9�r6�݌�~oA����l�SVͷqQ�#f��D���.H��#�8�>�����7��J��@}������O��H��y�O�y��Ffg���Gc���q؎�@ȓ�^rƩ���⠰������q���>�q�@��j�O"�3�TO�W��t�c�Z���ΚT,�:�J�ky{/,������T�&��� ̱ʲeJ�g�^IX��k{8ĳmo����~U,l��s*���C�Mv�<�lYXP����~�:�K���Z�΋h�Vw�i�����.h!�h�Z.k7�ӽ��s
��ԉZ�*�;r`�|Fx���N���4gA����H����]�`��!C��̢�`�$��i[��W�j�$��1��ENC�"_��Ü���xюa�����1�,��}r5�R�5`>`��H�����D�ۑ��ܻw�䑞"�[֪�vZcE0>F笰*���\֒y�P����ӻ� )ʲ� �L��|J�֑�&r�P�I������B�Gx�
w��ޅ��i�.��x9�v��A-r���t���_K�P�%�ȯ���P\m�ևu�X���i�|�C��.�d*�ɆUK^M���mC~3_;��^@���b5R��>Ų�pXou?�SD�p���X��gS�g�1�6��u��OvU��/��U6_����.����(����r_�Y{��w�w}jq*�g^��̄ld0�9�O?�;��c���ǡo�֯�'�#L���yϦ+U�L�,��W\g̓�����*��Q)�F�s�h4Ƕ��w1L(
�<���>����CX�4<R2"4�=(��=RF��%��gH�DԦ+�;LH�)�3T���%��|�0�(답:(}sW�����Hx���y3�f���}�!횦l�F��ҹNz�[�»Y4���F�mW�UȬ4l�G7�.OQ��6 q_I+����+���M!�����ܰ>��W�$�J�4"7j�t��WjoAv��շ|�Ȥ<�E�0�hVI>~��5�����;�@� f�CU8\4��0%8���;��A��d��%��\&#�G��!G���F�����L�zރR����w���>�}ΝRm�����َ�ѹp]�Gl�Ȧ�DbӨ���F~kY���.c}_1A*�K�
��6�|բO��;QN�"lzj���=��c�K&�g�ce�<�8�=�M/F�)b���+'���I��PW+���	���ZTNX[�:���$������Rcr� m�L���פzT��2���=�g��lZ�N��n'T�~�N�Q��w@�B���7Ȯ�N.|y	γ�#�]�T� ̵͌Ih��T�ޫr�[?p:p=�CF�^��Q��-s#�ڷ-��M����7��/�2${��G��Ϥ8��2Qp���W
� \�*Y��n	u_2���5!>=�Gb�Nv��p譾4�.�l*�lO�dl�z�d�Cz_o�"Xs�j�%Gs4���a=C$){՟l���O*���/%���dY�����~(t=��x���:2�K����x1ψȗ[��>��v�{׷ ��%mH�x0*�|$�伻���?+�yע����.$K�Z���r��G	/����^tG��9DyZ���F���׹�UP��^A��2�N�N�[A�/@C��l}9��X[�Gw���kD�C��<�+�Z��dړ�hmΆ'�`�w���z���?��� Ո��y�$4��=�?�@���5����c�yy#��]�[.;����d�W#4RKr ��S�!�j�C{��X�J����q��guʤ��� ~ �_,���Sb([�TW#���;eo�O�,�L����*;̭A�1��zUl�]���H�#Ϸ)?�2��W�s!Kt�M�Ȑ��K�¦71��vos-;B�
�@J��OA#7g2�.��DN	���;�o��7Gf�vr��骸c鎬 ��	�	pk_Bxh�08O�$z�pxq�����@��?��[���"����]���)�aP	[���dD1w�]j�|x�,�6��l��}�%�ӳ�L����Ȧ8{j�����=�Ȍ�1��z��T�Rhg�*��<�&��[��_�����3������FQ�4;^uX1�xZ6c��Z�0�`2 ��X�W=��z�^-�E�d�j���1͛�����W~����:l�!���eK��7+��@$!�>��V��*��i��a8�I����Ątm�;��Þ�W]nd��j�$��Z
�4��~S��;�<�k�f8��IÒ�mf(�Y�nJ _*+��RH�~���ZUS���,j-�d^������Te���������n�5� �G�i[��L0�\�����K��tZ��p�+_�݃ �R=���b���bLR��ǚ���1��R����N�Hx1�����������i�V�"��4i*S�����x,�<�1V�����|jv�ŜZ�gݨ�V:ew>̡.V�#�����A�b=�o�]ż���e�ګ��c\A]-�q��Qz��]
hu[�: ӢT��s�����`as �L���۩cU�T���)q�>�g&��:��(�1��E����,� Tzp��
��2�4p��k�����b����΅'T��S@=>�CY�fu���g��P�G�«hw�g
��d;�v�ˊ�(���9�����N��*9e}�L��甖m�� -`��n�{}ٰ]t6�
��=����
as���^�k�`�����>->9���DʬE;�l�>��ʕP#�L'Ϡ�r��Z�ި(m�(��ʯE���xϴn�u�1���~}O��o�����Ȏ4�V�%�8ռy�7�i�L�:mʁ�k��ri|���/��()P�A��V�^�	��I�D�L�����%JRL�lv�O�_����K���JMx
��%C}����!�~��QѹY��i������LF�i,cP���T>���K��7E޸V~!:������}5�_�~�?�'����d���dc��#��N��8wXa�W�{詇%�#*m���ğ�}�ګ	#Mqz����Ņj�9=��6_��.�Ӕ�tC6�^P��'�/�"������7n�[n�����0��uQ��jF?�?GNTxl��mɕ���#�MUJ��"D�+>�|u%��՚�E����0ג����3fKF�
��aF�_��DΔN�{�̡>�lC�����g�_woQ�k
�x�0�J9��v�����(��X{��)#��N��W��5$
tl��G��Q)¦����f�/�C�)�׳4���MyA���D(2�Du���O']�Fo�
I ��O�Q#��
k�5A3
�-���E��"	�n8�5�KTGM��
{��m!E=���ֵ�5�O����<r/ �O��uE]p�/��:&q*.�Da�#�j�x�è�L���R�_hϪ
`��*?���ܜ�4^4JhU$O��v��bVs:��j�'	fuż����1+X�9�x҄I���K�y��� �0#���DJ4�ҳf�]��??�⋉�6^��I)p̏���}�d(����L�γ���QԷ�d���<m��1�)˪6���M��*�+q�v&eY@��b4��Pn
�����N��%�K3dkUΘ�Q�����M���2C1Z�4$m�20f�tw�,U��~Ej����Z|Dţ`_�joO�����P�"�N��Kjӊ�sa3DI����p-��9���/h~��]=:�"��*�M
���+���"�r�s�F��`,�a�Lƺ%�!(m��dD?��L}$3��.�͊*ˤK��8C5�oܯ�sY�h�g�&n?��< �'�{t*�4;E��\1��9i!Ȼ���P2����j�P>Ah��$��v���Y��z)g�����99��2ui�"B	\�S���<�{
K�o�����I�r��z�ߑ��\��m���w=�ҋ���B9Ѽ�|e�"���3~��>q�őA1�H�������%���ɗ�*;9���w�wb��1��Ka���2�q�lc�p��|�~������R�f�U�6�}�U����y����,Ni2T�
k��xAG��D�Z�Q&ɃkLk�h�M�Pճ Ν�[�&�@�'Zf
XlxV65EB    d975    2580��l���e��E�:�K̨���̤�������O�?+I��s���j���5�A�5�T� F����Sj9�|C����͂��z���tO��"�+׭��������E3��ڱ�9]�z�;;cwV/��I�����2��s��G�׉朆��v[Q���č���[hU��r+�� {��ӇM�*����+� ����*f�J�s�?L���l��JzJ]㳶���Jh�vW�+m-'�x<��o�=�k�M����X��w=���x�S�$�������J*��'���%ҞC���_�۔�ȍ�u�+�d7ujʃC$�V���h����u��	
�l�u/����ג0�X�S�Lx����e�4�_s-\�C�)�Z����f����`����2��sJi%*���۳�J;V?g����tA�C�&�+a��vX���s�����1>pr�',0�_^��B9fa�qа��rVBS?�6p� -�����QzJTW�vbP�; E����݅����0��v�����h����!��5p/~'˾���ԉ�.��,B�:��XAx~Nw�[eľ�m��΋q�K�0���[r鎖w괔�&�D�ֺ�K�>����"C�P\S}��jytPM�#{� ��;���u]��#Ӕ�g���$ L��p#��+����u4���fS�@�ԳG�����I�����$n<s�K5D��X���u��j��Q�Nd'5i� X�q��µ*�D�T/1���f� ����h�U]���~�]�d�P2��٪b�	��,f������1�yC�1u�a��T�X���ht�C��G� I	ը.)#�mًP[��"�$�Oz��w�#�����!����I'��R��y���A�'��1�b��e�0�bx�
�O��k9VmP��^�D�@+�gZ�0��b9磉^��� 6*)��x
���}Р�H�V?�:�?��[�r��? wi�y��b��^̕�D����4CI@ۤ���g��s�1:��{�J���B����ɱfO����+�x���]���/�?8<��!Nt$OS����	�����
�ޡ�+��}ɴ�5��p	�0K�����0�ݭV���7t���v�%r������P^A=�շ���`��?D]y�[��t�����E6�Ss7PGV`�4����W&URu%���!NÚ�$�B]�?}��g{3��h6�=G�JH�F_[w��rR_���=�?�!>����Ca��>܊ڣh.��+dV�9�&η5��構К��H!�����~����E���#�׎���+tqR�8��8� ���P�.��A�P�օ��^�H7��2m_�kKT�ʰRuG����s|�G����~�"i�ԓE�0]�t-:�DTy������f͘_���W�+|1RG����sݷ�(Tx/�d��Z'!�s�����t�dn.Ҡ�I�i}����]̄�d���~���U���sf��fԧ�c;hë��N<Z���bP	�Aq���N���=�$��;O8���(z����طH��I����<H �8ǆK����lE2]ƻ�j�������N�_cj��
vg��p���r���\i�ؑ���U��Z�%���4É�膯�Cg�������C��z,�I����|Y�َd�FT��R�zRmq�s&��f�	���{�yŴK��t��?�儾E#��@Uw�̒ 5�����|6�k�fj�is��q?�hS5�N���/\d�+�8��zJ�+X��D�O�����R7���:�����Im�%zZ��Z�>���Ɍ�x��򽼳C��`/�*�����̨[Qf4�p;�;:!�M�D�#���^�\L�s�ܭ����*nҭ��y�yئ�����*�
US��l��H���$!�@Q�M��=�'�*Y$��x�%�R��:��l�6��Bn����/��LT�%7N���1�s�wFi�.fE���[OՇyP���`6�(�ϧDW����,:���8�Xv�^�%d5̙���S���Eς���cX5��_j�lYdq��Xd�EB�ԟh꼌��1��B%�m��=���ҏ�K� [��2Ybl�|x�����K��S�ܧ,IK�nE��j�,��elLL��Lȧ�7���S��4�k?�-��h�Xe��U4�M �1(��UT܅j�`A�8�;�K��s�VG`�-������u�)�V��m��يR]��T����?��p��[�� p�C�!<�6#v�}��_/[T���A��5d��]`OC%/A[T��jIϡ5��b��3�^4�"'��	��  w�����G�4��J���2��cBa`���	�MH��WR>��t}��+	�_W2�}�XJ�[��8U�ma������T��Q�<UXb������Q�i�i=7�]�"|N���%CГ�#a>6��/�i���>*b���^�Uo�y�G�L��m@p0�1���~���M�5�5�;���i~���H��]Ψ1��Y�41��UU�O��Y  ���S���M�)��o��8��W�0���!�l�"o��{��ݗ ���[[,T��!ȅ����W���ޔ�ڮh:���H�4�6M6���?de�|��۩k�!mͷqTI�y0=`**@al�8 l��j}�>!Ă$��t�R��z͍�8��6��k��bK!PĿK%����x�y�V&aV�9�(��8��9&7�ڵ��K��_́���4��#���A��ڿ]���9����#` ��>�Iv
B�{�_aU�J�ea~��6y�T۪�	�u���nS�v�0�ۿR4�w[�?�U�9N����D
�L>�B23�e/z)�+�
�?jq��4SM?~0t��^�7��*5��1���	�#�b�K1�_EZy�#��r��Io
輦i�]�� @��#F ��U �V�T��������&$��X���[�^����@Ym�Ά�Zz��)��7� �y�2=�3�o~�b�q!$��$�Z �����SCw�Ue��(���Ws�k��V���*��zI��hE+ȽF�D�mp�������G��A����R:��<G;Tż��"g�AA?\��4�B5]�1���s�k�,��o� �Y��D�Օ�y3<���!������f2,�e}6��{O�����C�U5�z��m�_�3H1ܻ��7�t����`��8��3�p.�= ���l�>{h�ʉ�	�Kd��]*�y�!6B�:I�ěN�r�\��3V�ӧ�W�g��o��7�Pu�����Z_�S|�W�9���9�|��q�I�_>��5�mꙟ���F��m&�q'�@Ӎ�!�3��z�5~���H��:��^��%m��0���7�0P�ţZq(����V@����W��.
ʙ2�U�$�� �#= GM���@����!�9����I�mh���5ݍ�����q�9+�(��og��[3��5���ž>Y�n29I�!��׭�[ڔ�5MF����מ�� p�k"I89�_Y���M��`Ҹn�ꑢ_��s�k �����������?����Ʒ'J��)�W�}�>x+��;.� Vo��� �<?8�Y)MD;� ��.ĕ��S,��[����̎j���L �!0aAiOڇ��N"��ߵ�C�f���UkE����`顄yd� t���N#�{����o/iG�ktDpy�@��>/��'z�A�4H���AFg���"���,m��[D� ��d�"u�c:���>	 ��� ?�/����[8��}h+na���y�L����R�qW��9�����=����r6���<L��-�UG��ʟ�k�sC/sP����dI:0��-�/t0S�#n:�8�%M)���b�!�q7��d$��d�Q):E�Ȏ�B3VЀ�>;�K�ћ4@r���C�'_%�4���{� y�Ώ�e�r(0nb�'E-e了��q��R��ED���	�?*�`�"�h��k�ރ�UF��-_�Pؐ+�У�����j�HRu~�R&=\�ަ��ȯ[6<��m
$z^M���JUgV-�7��R���~�8��%��wS���@V�}��m��T�ٰ}��9Ĵ�F��Ilp��T�����M���hS�T�/�H�~�M���#�W��9,<8�-�VC^��L�l4��w��T%J�#&��bi��bCUq(Jy�㷐�Gq�a�@����r�旐�wx���C�`�jzen�\j_�R]��h�_^���7�/��H��Z�hr}+1�G��q��Mm9��u�l�:	�6k�b2\�P��B�c��nE��.�����i!8��̦���Z/�uF@j��?���W��8���
�mnP��E���O�[P�Wu�韦A�c�dp�j�C;�
�v�R��P������%��� =�$� \��k�&g��F�����Ԟ�|�qi�Ql�b���5\�<�Ka�N�b�؞<��xbcy��������f��M��o4?�)~=$A��gQw��Mu���y��"�4�T�����ӓ���V�\�W��>{DTn�v��+�jW�ɫ  �Ńj��[pu� M��+����b������u<;�Y5j�w<rn� ���O7K�f�z#�+�� ���}q�_�Ğ����W�Dׯ��q/��M��
X�~	أ@�Y�w���ʺܯ_ti{8�tmM~��k�&�W�
53�,����c�����S7��l��������p��Z����>�B)+�[:���w��Լ��b��������߶G4K [c��`���iPo"���@�}83qq'b;�Q���κO�1-m`}9i�kڎHd�..}�-�v*�i��)�U�|T�����D=� g0�=W��`o�6�g�a����΅2���z�"�+�]	�A����X&
�8;a���v���=��Թ\����G�#ikbfr��DR�>.k�HѢb^`G�M')�(8w6F��qW��r<4�f���)(��mX��A j���x�D�����gfZ�	����>����S����i��H�ő�J�I{R��RN���
���K��۰}��B3���݊I�c���o�-~���
Z�a���w����k�?�&�$Q���� H�K��E9�f,N�@%2/�� ���y��&�e�����<����:���b 'R�
3ך�5���]]{d��\����FV4Ȥ#Ǽ#2�#]s!��L��j
�Xl��?*'��1f�p�u�X�d���G�;b��cT�j֡=�O���R�/�1��7�����W\`;���s(���,<+we�B3s�e�B���'ʃ����`�J5b��_!oF�_Ԋ����6�`wYTC��_:�bNץjBaR�f#�i��@�nvω"���jR��衙��w�$
,?��Br�ܻ�=w)��8���Ux��=�+�kڙ�I���Ď�p�4��A�J��O�x;��>\��XD�����߬������Uq �;Q�Pz	tV�R�͌R���h�Wc���K�5W�����F�Lh�����/�3[��.>�}�}�>l]ǧ�L�O[Yj�L=Uz{�8ƈ��c���.�;��rDM��?�k�S�d�v.�Y�p�2�(F�ƚ=��'��ޯ�&fryKw�Lރ�H3��7lXG��z���Lu���+`'L=�Jw�m�ۊ�RB�ܪ7D �6�! y�`���	e�P��H��wCZ!?޸��q�[)�}?R=4�r \wp3��#�+�y��s�JY�ĸ?V<�4�mX�5v|WKU�"�y6�m0�����������,�k����H�J�+�H���h�cQ!�N�!�F-�W :������hIL�{��.P6����֞��V���I�4;����!����H��5�#����]QP���ߟqdMu�����<�爔j!�b�J4������N�e��!�(����)p�����́�[GaF�͈h"3�	1���E������$GM޲Xpʂ�Y��m�.�+�yY�!V����#��f�(�����g��X�Q^���)���[t�n��i �1Z�-�?�A�q�pF"
���?U֖s�'>�~'eJ��mJ�����ڿC{ƾ������.��?��={��-�����F���[�	;�4��|=^�I';3��2��Wmy[��m��T����݃6��;ӓN���z�FX�"Gp��O��[�D�\�O釪�dd�[����'?7$���R�%zP˂�#$!�O��;��q�Y�w���j+��U�2�!��Z+�ut�	7�����VD8�}�F�[׍�����T�i#�<G�?�x�Kz����������N] �U:�ɮ����q�"?�cV&�$lYe�\���4$��vd�2�>*6��̧�ׄ5xg,�Wg��)�P�՚f3���Q���Oɖ��%re},��`|��Uv_]n���������&��d��W����D�����^�f����r����Ĝ��J�ņLJ��E5@,Z*�?���n�3 �˽C$��gst%1�/��4����Z�"�^�*��M�<�Jc��)����.?���2�$�\��Ց� ���g�~C#���@Β��)��TJ1��B观�@i�f�����2�g~,�`��eEjW{P͓�䂴k���A\����U�L��3l�a�|9\�$�"|��l�%M��ϰc ų4$����������ɿ�D�\'��6�or-�����$9��)�G���c ��Ų�R��6=-�����q�=�p��=k��(�D�hn�v^�P{��VֵŬ�˼��6rZ�~07���j=l�� �2tլ��ɘr?u�	r�r^8�
����C��]�Xr���|D�E�����ײWν�ڒ�[9c)˿���N�va���+r,��A����:���w�-�4xgZ�U�ؽ�5.K�{�yKQ�������>?1E9h����w����ф�<i�K��	f��Kx�и�QS��;ڲ�lc�G���U�7��p��fY��><J�R�ts���;��EL�77�����.�9M�@�,sa 8_d�=���+�p���$���ƍ}/���o��)�'J�}����/�,�eX,�j��Q����Q��ڥ�N��Z�&�E���+:�l��Ξ�؁�� z_D���?�%���`�4��,lK����ֺ�c0$�7���C�	�+���Z)w;9c,�ٸ�\y�l_1�'��+F��N��n1��NW꿭����Ѓ�Ȍ���8�ث��[_��&ϳ�M��>9���B�K�*�d�BB�/w�%�:��$J�����K���#f�>I�K+aD���?R牅�e6g.���k��� ��OƏ�����?��rOǎ�Qr�7�n��Ρ��Q^^IYx9�	�%����(�hմa��2��E����ݹ�� ����>���������^�MYJ����~p�b�p������i���ڥ�r�V����n���-��p{�<�D�8��h�Oڱ"��d7��:�˽_KY�2+�Py��_a�Ȟ��F���W���k즎��D�1QOO��x��;�����?ބ�á&�����w�H�(5���)�W־���_�#s�c�L��B��>�B����,x����&1ȋ�C7���,��,H��Q���Ȗ�*W�����b�h���`jw4��-K/e�m�}�)pVr��1�A�u���A��N��n&-:x>gU�q�I�ل@X����ɣ�5['ހ�<M��u���M�n� K�I�-�W�H�L�����u�8�5�<-�s)8b�$�x;���D̮鿭�W��x�7���~��7�(E�}A=z9�7��;@Ɇ��t]�c��T�4�L
^��m��N�E�=�P�4`�0*��$(�	�kE�-#�:�f�)E�UYbL1Es���l�O.#����g�Ҏ(9���%���H����(Ѱ�3LAv��{+��⨆�9e20��.Ja�e�&)���$^]�tډ��̊3dc�k(?nv�I� ��{��e&X��\���R_��A��%�W�=f�#�|�.F= ,���xj�U;�	w�G	��K�k��n��;��d���
q���8d(�s��g���Hj�8aע5B����i�C X�zP��F%�����H����ړķJD?�����]�{��\�2\�m/��n�ޚ����_~���Ai�/����N��c�g����}���0� ��΅�9�t�����S	3��!��5�h.�x�Q9�p�	Ɉ+1�8"���[���i��{G�3����"�~	������ܰʬ~B�=���'�bf���]|!��0gZ���2�\�!��"MAg�������Ū�6혈 1�+`l���~��ק���]�^0A��=�0�w�EV�L�[�����8�8��T��9ѵ?H����kk�X���8���O�I���G[�bp�;���/�ЎV�'\��k�/��Yi��Z��8�1�Y�*Y>/�>t��Jj�iJ�o�C����Ȏ�8k +E���GA��x�GQ�����}��1�pԦ;�+����o�v�J�P�M�ܻ��S7� wu�Y��/�܆��L/(�ަxL"���Ͱ8A�\�����볰aj�XӑB������EJ:�'n�r&� �FT�����i�1��O��=�A�����9�5H2)jE�(^�آ���w-n��H0 ֡��AӪ�c3����tP=�ц���k_w�,g��w��ܚ�`�#[l���Ӱ�M���Rf_3��"���Q·�
���0^'O��ө��*�f#���k�9ݠ�v��� �X­�Қ�/��\~��0�Ȩ���~^���i4�i��v7|�BIE�.� 	�DL9_����Ve��R�	y�H`�[d,W�w���6��l�he_�lcH�߫�n�W�}���eQ=��M�hzGQ�Q���o�=g�y&�����Ŵ���m�(��"��@������?�*�r�y9�x�i� �ر�4��:疜�3�8Yz�?̷�����b������wM0���&?�,X4�.�CF]eȆ�}�c.�OX#	eh��A{� ��)��#lƕ�L��hg�>sxX�Ob���e����ỉ����N�����r��w� ��rZ�4)"���U����%ד)1PR��q��j�=C�I^��r����#�=LF�Ĝ��Ԟ�	�-�+� ���p� �����M�nH�c�=�L�0Oc���8���c��s�Z4����=F;������FMV�7� >K�O��?�,�oI��$��Ш':쓶���Y5?�P|��{����èf
���⠀�ނ
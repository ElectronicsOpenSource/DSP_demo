XlxV65EB    1e0a     a00��/#��wk��\�D�z��P�2Ɩy�Q�~�W�qʙ}�2�z)����W&��wa�F�9 Èʈ�pTF����)	@2Q����Vw�[����C�:2ǩv����b]�i\�3�V���j�^���g>10w����`#��@b�	h.$�k�H�H�?�F�hXd�-��pH�y��M�B�5w�õ�8���ݿCb�j緮�ȫ�ds�
����#l=3�-�?�6v�N3� ��?�ݜ7�;p?�k㙗;�X��/@S�Q�#9Z����&$7^WB�ɹIaf 2�.���*Q�r�N�B�sχ
�_�c�����WVMOEfm1�#LS��ǟ6ȇyP��g��>�Ln��,�z�h�}�U��h����V�0[ݮMxT���WE���gxHS��X��x�����a���<O��B&����=��0��G(ķrY[�l:��4�� ��̹!9�RT�6���mV���ӯ��
v<
��c�1�9���(�ʹ�$����i��tC�5s�a+�$�X;�o�z��!��wJ��*]�w��=Z��}�o�͞0��_�Y_�r.�G-l�����y�@���h�����V���$�3�ǩ��{}�Y��0s���t�t�^�L������X$���:���J*V̤��'PX-���Ξ���s�ꌁj�HAo�������+uע�`��O�F�� ��&�Q�'�NQ�]���|���%�p�F�� $V3�lm�\W~�HH��Z�	�vu)�3|,�m��P��,�9�̌ق3�"O/;I�8���vDy�[_�\�u=����81�V��ަ��xޏ�W��J��i�Fw��!Iq�{d��y/tx�>����mD�����o��Z��*Q)I�8��9��O���(�����ʤ=�\����]8H�,y��-��1�}rI-�L�ki�&¤������B)1���199� zܶ�_i7 �^�T��㌺2S���E��%�$Z5�a����J���<eo+?�%QY,�V �ڟB�k����!p��x����3��� ?q͍�0)������>�8A>B��yN��/�~tM�\{�t��B�j��� �V���[s!5}4�\���d�=�eB�Sb�kHj����?B�c�7�'⥑��^�����,�W?�����-�H�,˔��ܔTU�s���+dD�Ռf���½�~�W�>����{��Ɂ�"�M���b�a�;�����=�O:��ud�L�)Q�g�l ���r�����W��ޮx$h�g�]�I���[�T���.� ��E���tuB�F���^�0��?��?�� �ok���)G
g��{AM?��M>�kؐ�Ա��"l ���_�o�Z�{�&��$/�����8���p�'ߤIނ#��RT�ڪ�� ���?�c�o;i���Ȉ��Z�_V	ЇәN�E0}0��g*������WH������D�r�t��-	if*u�s�BN�e���	pJ LI]�2d$9��z?�玬
X���u�ޥ���X���o�u@��n1*�s�B�g�1�^�}n��ƐZx[�Z7$�O���h[m���/9��g��o�SY����p�gM�Օ2��9 y�(�H�tE$��K��b� $4����k��r�9���u.��߇P��i'�����+u3+�ew�X�3f:��)��`�u|�����茵#�A��p��|�Ak�!��Yߘ��C༣YaJ(k���i9�Ϝ�Լt+�"����*r�p�e3�k��AL�Q�;k�/7���WB�[C6��楹�n�q�
%�V���R_��G� ���H�����?F���3��BX�U6RL��6�}��"&S��P�u���1����>j��߷\B8N�����<��CP�q��p��*#�UM�ʖ�a�ڌ��L�mR)L��[t��`=}O����֕oY���9��L{�F��C�ٵc8�űܱ�O\�q�`�׈�(1/nG���?�6���ܘ�2ܞE1yd)�~$'�pV�[B��F����W�0��M�A�C�J��P�#k�}�o����M�ZsU�c*h��H�e�PG��.����D�b��l6mY�!оՎ7�6��əp7�����Ŧ��*��z/<L�[������.ع����_�`t��D�^�>��;F�N��-*�t���3��8G�#T�R��6�wAY�R�V\�����z���?l�5Q��M#K"D;լϕ9�I�,S~�_���Sr�͛������6��=��OCB��>�ҿ"�8{2,Xe��N��նy7!Q<���÷%�ȦjN���[�0��4�1����ʐ�D?�=�!�Ӻz�sn�g<1;IIIR���;�r��hO ���yS��k�@s��5�Q�_�;���F��S舞E\�Wj�?0��|d'g�*L?M7h�WdC�`;���e������t����?��9��C�x:�̧ߌC:�Z�$|m��Q�4����ZEM��]�*�\r^Kzi+оӆ@�tFD
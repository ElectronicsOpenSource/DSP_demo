XlxV65EB    31c0     860���[���@��$uw�l��w�ׇ����L���S7��5�R[-\���\"�%2�[n�(1��]ҽ[\V
�o��R�=z��Z�X�V��H�˃����������w�x��߸38"�s�c�	��^��&7�z:E��e^�*'g*)���ށ�"y�Y:����M������s�����2<���!��}�4�"i�d-��}b�"[;;?ir��Hő	t#d�Mz��g���C��@,���U��V�����Y��w��$��t���ƺ��5��X�(��~̽���;�w*k/Ikb���`���Q!"Sr5�+����ˊ��N\�o	*�W�S��2z>�)B�hܟ{\cq�)
"�|�� ��6Sb�	��"
�!.�QD�s�\$��s����ke�z�6/6�y�	��<��U�����m(W�!a��7ȡM���Ӳ���w�8�m]� s8&�Y��U�0R��W�z� D�44@3���N_$#vYt,HE�����-�������b��W���:������FW���O�'cq�����n��R�߬r��.]������H�I'�Z��8&�=T���]T��!�ᶺ/�Xz�)�	~x~�����o�~Cm��Q)���~e�ɫӆ7̅�CK�ӆ�VFi�=��'���E�@��tݕ�(�^���VA>���N�E��09����_E�3%y�O�5�#r#Cv�ϷN�������J_!^w8e���;h.����;EVS�PP'$�#w7��S��%�������9]��7��2-u�'�LG�-���/��H��k���x�y���k�>R9B/�[Q��P���WYŽ:����A��\jÐJ:�H�Z�&�f7��h��mJ�?\cs�.���ܓ9
�}Z+]���̇�	2p��=�����"��$��N���U�hl��-2�dY�0��(t&�1�k�����c��%�N���u�+��"��0��i7r������5WiS_��G��gZ�k`����e5Ҁ� ���0�#�Qe�4�����|�6|Z�#cJ���OB��K�̌K�i*D�P���ud�y�c�����14q�z��=·��<��2��U�(Cl�$;����Y�|��yMg#��S�s�{�.�UJ���o�s�O�P}a�������`�5��S�U_)6��c���C"�o����l嗸d:�k�i��z%&�}�a))�&�e�C���䀩�0����0�#fr3�pH�u�S��"����!_`2�{T���!X�/IO�.C�-���Qz��)�g�������J�'g���y/RqR6�}`1O�R��T����0�Q��[�â%ȼ�L��$��I�V`P�ئĩ��d��M�`�����<MH�<+��uѬ�<�5|�����bW�9�"'[��(K�4�(aT�*Pg��7�@�N����a�E_w@���t7^�����;����]6�ѥ�S+�F�勉�/��,u0q�4�mf �\����m}�D-�GG"�$�$�Wq�d��6��}	�����Dk�.�хy��P����"y�X�<E^vi�U4�.����� A���}��@H�B�]��9T�9��y:�N}Kq��]��u9~xv���A)<�`�x�{�8O�m�4�Q�d{w��ƿ�=5#z'����1��*�OK���y�6ˁa��?��3�#|�)b�(��ì�F:Ѻ,j�xM�}�2� /6�m9���H����^P�GyJ�w^���5H/��G�S! ��$�6x�8�);k^�l�y�eN*Cߠ��ȕ?S����+'Z�m��rc��Zub #���g��������l4�&���a�^u{��'"�Thm8`ɵI���x��}��w7v/=�������0v͡� ժF�3:V��`M��l�[s,��˭ ��@�d���d0�ի�S����x����)dH�T)����M�`Mj��R,.	@�R�]����l%�m�	�vq}�V4AeZ��ֹ���!ѯd�#��]�˴�db�*��֦}9YP�alV�?_z�������6w���"��	��	ߩ#�^�hr�c�ޙV�V�PA��p��1�9�}JBp����`Q